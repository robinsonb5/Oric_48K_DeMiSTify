library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"7f7f3018",
     1 => x"36634100",
     2 => x"63361c1c",
     3 => x"06030141",
     4 => x"03067c7c",
     5 => x"59716101",
     6 => x"4143474d",
     7 => x"7f000000",
     8 => x"0041417f",
     9 => x"06030100",
    10 => x"6030180c",
    11 => x"41000040",
    12 => x"007f7f41",
    13 => x"060c0800",
    14 => x"080c0603",
    15 => x"80808000",
    16 => x"80808080",
    17 => x"00000000",
    18 => x"00040703",
    19 => x"74200000",
    20 => x"787c5454",
    21 => x"7f7f0000",
    22 => x"387c4444",
    23 => x"7c380000",
    24 => x"00444444",
    25 => x"7c380000",
    26 => x"7f7f4444",
    27 => x"7c380000",
    28 => x"185c5454",
    29 => x"7e040000",
    30 => x"0005057f",
    31 => x"bc180000",
    32 => x"7cfca4a4",
    33 => x"7f7f0000",
    34 => x"787c0404",
    35 => x"00000000",
    36 => x"00407d3d",
    37 => x"80800000",
    38 => x"007dfd80",
    39 => x"7f7f0000",
    40 => x"446c3810",
    41 => x"00000000",
    42 => x"00407f3f",
    43 => x"0c7c7c00",
    44 => x"787c0c18",
    45 => x"7c7c0000",
    46 => x"787c0404",
    47 => x"7c380000",
    48 => x"387c4444",
    49 => x"fcfc0000",
    50 => x"183c2424",
    51 => x"3c180000",
    52 => x"fcfc2424",
    53 => x"7c7c0000",
    54 => x"080c0404",
    55 => x"5c480000",
    56 => x"20745454",
    57 => x"3f040000",
    58 => x"0044447f",
    59 => x"7c3c0000",
    60 => x"7c7c4040",
    61 => x"3c1c0000",
    62 => x"1c3c6060",
    63 => x"607c3c00",
    64 => x"3c7c6030",
    65 => x"386c4400",
    66 => x"446c3810",
    67 => x"bc1c0000",
    68 => x"1c3c60e0",
    69 => x"64440000",
    70 => x"444c5c74",
    71 => x"08080000",
    72 => x"4141773e",
    73 => x"00000000",
    74 => x"00007f7f",
    75 => x"41410000",
    76 => x"08083e77",
    77 => x"01010200",
    78 => x"01020203",
    79 => x"7f7f7f00",
    80 => x"7f7f7f7f",
    81 => x"1c080800",
    82 => x"7f3e3e1c",
    83 => x"3e7f7f7f",
    84 => x"081c1c3e",
    85 => x"18100008",
    86 => x"10187c7c",
    87 => x"30100000",
    88 => x"10307c7c",
    89 => x"60301000",
    90 => x"061e7860",
    91 => x"3c664200",
    92 => x"42663c18",
    93 => x"6a387800",
    94 => x"386cc6c2",
    95 => x"00006000",
    96 => x"60000060",
    97 => x"5b5e0e00",
    98 => x"1e0e5d5c",
    99 => x"c9c34c71",
   100 => x"c04dbfe2",
   101 => x"741ec04b",
   102 => x"87c702ab",
   103 => x"c048a6c4",
   104 => x"c487c578",
   105 => x"78c148a6",
   106 => x"731e66c4",
   107 => x"87dfee49",
   108 => x"e0c086c8",
   109 => x"87efef49",
   110 => x"6a4aa5c4",
   111 => x"87f0f049",
   112 => x"cb87c6f1",
   113 => x"c883c185",
   114 => x"ff04abb7",
   115 => x"262687c7",
   116 => x"264c264d",
   117 => x"1e4f264b",
   118 => x"c9c34a71",
   119 => x"c9c35ae6",
   120 => x"78c748e6",
   121 => x"87ddfe49",
   122 => x"731e4f26",
   123 => x"c04a711e",
   124 => x"d303aab7",
   125 => x"f8d7c287",
   126 => x"87c405bf",
   127 => x"87c24bc1",
   128 => x"d7c24bc0",
   129 => x"87c45bfc",
   130 => x"5afcd7c2",
   131 => x"bff8d7c2",
   132 => x"c19ac14a",
   133 => x"ec49a2c0",
   134 => x"d7c287e8",
   135 => x"c249bfe0",
   136 => x"b1bff8d7",
   137 => x"787148fc",
   138 => x"1e87e8fe",
   139 => x"66c44a71",
   140 => x"e949721e",
   141 => x"262687f6",
   142 => x"d7c21e4f",
   143 => x"c049bff8",
   144 => x"c387d7e9",
   145 => x"e848dac9",
   146 => x"c9c378bf",
   147 => x"bfec48d6",
   148 => x"dac9c378",
   149 => x"c3494abf",
   150 => x"b7c899ff",
   151 => x"7148722a",
   152 => x"e2c9c3b0",
   153 => x"0e4f2658",
   154 => x"5d5c5b5e",
   155 => x"ff4b710e",
   156 => x"c9c387c7",
   157 => x"50c048d5",
   158 => x"f5e54973",
   159 => x"4c497087",
   160 => x"eecb9cc2",
   161 => x"87f8cd49",
   162 => x"c34d4970",
   163 => x"bf97d5c9",
   164 => x"87e2c105",
   165 => x"c34966d0",
   166 => x"99bfdec9",
   167 => x"d487d605",
   168 => x"c9c34966",
   169 => x"0599bfd6",
   170 => x"497387cb",
   171 => x"7087c3e5",
   172 => x"c1c10298",
   173 => x"fd4cc187",
   174 => x"497587ff",
   175 => x"7087cdcd",
   176 => x"87c60298",
   177 => x"48d5c9c3",
   178 => x"c9c350c1",
   179 => x"05bf97d5",
   180 => x"c387e3c0",
   181 => x"49bfdec9",
   182 => x"059966d0",
   183 => x"c387d6ff",
   184 => x"49bfd6c9",
   185 => x"059966d4",
   186 => x"7387caff",
   187 => x"87c2e449",
   188 => x"fe059870",
   189 => x"487487ff",
   190 => x"0e87d4fb",
   191 => x"5d5c5b5e",
   192 => x"c086f80e",
   193 => x"bfec4c4d",
   194 => x"48a6c47e",
   195 => x"bfe2c9c3",
   196 => x"1e1ec078",
   197 => x"fd49f7c1",
   198 => x"86c887cd",
   199 => x"c0029870",
   200 => x"d7c287f3",
   201 => x"c405bfe0",
   202 => x"c27ec187",
   203 => x"c27ec087",
   204 => x"6e48e0d7",
   205 => x"1efcca78",
   206 => x"c90266c4",
   207 => x"48a6c487",
   208 => x"78f7d5c2",
   209 => x"a6c487c7",
   210 => x"c2d6c248",
   211 => x"4966c478",
   212 => x"c487fbc8",
   213 => x"c01ec186",
   214 => x"fc49c71e",
   215 => x"86c887c9",
   216 => x"cd029870",
   217 => x"fa49ff87",
   218 => x"dac187c0",
   219 => x"87c2e249",
   220 => x"c9c34dc1",
   221 => x"02bf97d5",
   222 => x"f4d687c3",
   223 => x"dac9c387",
   224 => x"d7c24bbf",
   225 => x"c105bff8",
   226 => x"d7c287e1",
   227 => x"c002bfe0",
   228 => x"a6c487f0",
   229 => x"c0c0c848",
   230 => x"e4d7c278",
   231 => x"bf976e7e",
   232 => x"c1486e49",
   233 => x"717e7080",
   234 => x"7087c7e1",
   235 => x"87c30298",
   236 => x"c4b366c4",
   237 => x"b7c14866",
   238 => x"58a6c828",
   239 => x"ff059870",
   240 => x"fdc387db",
   241 => x"87eae049",
   242 => x"e049fac3",
   243 => x"497387e4",
   244 => x"7199ffc3",
   245 => x"f949c01e",
   246 => x"497387d1",
   247 => x"7129b7c8",
   248 => x"f949c11e",
   249 => x"86c887c5",
   250 => x"c387c7c6",
   251 => x"4bbfdec9",
   252 => x"87df029b",
   253 => x"bff4d7c2",
   254 => x"87d0c849",
   255 => x"c0059870",
   256 => x"4bc087c4",
   257 => x"e0c287d3",
   258 => x"87f4c749",
   259 => x"58f8d7c2",
   260 => x"c287c6c0",
   261 => x"c048f4d7",
   262 => x"c2497378",
   263 => x"cfc00599",
   264 => x"49ebc387",
   265 => x"87cadfff",
   266 => x"99c24970",
   267 => x"87c2c002",
   268 => x"49734cfb",
   269 => x"c00599c1",
   270 => x"f4c387cf",
   271 => x"f1deff49",
   272 => x"c2497087",
   273 => x"c2c00299",
   274 => x"734cfa87",
   275 => x"0599c849",
   276 => x"c387cfc0",
   277 => x"deff49f5",
   278 => x"497087d8",
   279 => x"c00299c2",
   280 => x"c9c387d6",
   281 => x"c002bfe6",
   282 => x"c14887ca",
   283 => x"eac9c388",
   284 => x"87c2c058",
   285 => x"4dc14cff",
   286 => x"99c44973",
   287 => x"87cfc005",
   288 => x"ff49f2c3",
   289 => x"7087ebdd",
   290 => x"0299c249",
   291 => x"c387dcc0",
   292 => x"7ebfe6c9",
   293 => x"a8b7c748",
   294 => x"87cbc003",
   295 => x"80c1486e",
   296 => x"58eac9c3",
   297 => x"fe87c2c0",
   298 => x"c34dc14c",
   299 => x"ddff49fd",
   300 => x"497087c0",
   301 => x"c00299c2",
   302 => x"c9c387d5",
   303 => x"c002bfe6",
   304 => x"c9c387c9",
   305 => x"78c048e6",
   306 => x"fd87c2c0",
   307 => x"c34dc14c",
   308 => x"dcff49fa",
   309 => x"497087dc",
   310 => x"c00299c2",
   311 => x"c9c387d9",
   312 => x"c748bfe6",
   313 => x"c003a8b7",
   314 => x"c9c387c9",
   315 => x"78c748e6",
   316 => x"fc87c2c0",
   317 => x"c04dc14c",
   318 => x"c003acb7",
   319 => x"66c487d5",
   320 => x"80d8c148",
   321 => x"bf6e7e70",
   322 => x"87c7c002",
   323 => x"744bbf6e",
   324 => x"c00f7349",
   325 => x"1ef0c31e",
   326 => x"f549dac1",
   327 => x"86c887c9",
   328 => x"c0029870",
   329 => x"c9c387d9",
   330 => x"6e7ebfe6",
   331 => x"c491cb49",
   332 => x"82714a66",
   333 => x"c6c0026a",
   334 => x"6e4b6a87",
   335 => x"750f7349",
   336 => x"c8c0029d",
   337 => x"e6c9c387",
   338 => x"f8f049bf",
   339 => x"fcd7c287",
   340 => x"ddc002bf",
   341 => x"f3c24987",
   342 => x"02987087",
   343 => x"c387d3c0",
   344 => x"49bfe6c9",
   345 => x"c087def0",
   346 => x"87fef149",
   347 => x"48fcd7c2",
   348 => x"8ef878c0",
   349 => x"4a87d8f1",
   350 => x"656b796f",
   351 => x"6f207379",
   352 => x"6f4a006e",
   353 => x"79656b79",
   354 => x"666f2073",
   355 => x"5e0e0066",
   356 => x"0e5d5c5b",
   357 => x"c34c711e",
   358 => x"49bfe2c9",
   359 => x"4da1cdc1",
   360 => x"6981d1c1",
   361 => x"029c747e",
   362 => x"a5c487cf",
   363 => x"c37b744b",
   364 => x"49bfe2c9",
   365 => x"6e87e0f0",
   366 => x"059c747b",
   367 => x"4bc087c4",
   368 => x"4bc187c2",
   369 => x"e1f04973",
   370 => x"0266d487",
   371 => x"c04987c8",
   372 => x"4a7087ee",
   373 => x"4ac087c2",
   374 => x"5ac0d8c2",
   375 => x"87efef26",
   376 => x"00000000",
   377 => x"14111258",
   378 => x"231c1b1d",
   379 => x"9491595a",
   380 => x"f4ebf2f5",
   381 => x"00000000",
   382 => x"00000000",
   383 => x"00000000",
   384 => x"ff4a711e",
   385 => x"7249bfc8",
   386 => x"4f2648a1",
   387 => x"bfc8ff1e",
   388 => x"c0c0fe89",
   389 => x"a9c0c0c0",
   390 => x"c087c401",
   391 => x"c187c24a",
   392 => x"2648724a",
   393 => x"5b5e0e4f",
   394 => x"710e5d5c",
   395 => x"4cd4ff4b",
   396 => x"c04866d0",
   397 => x"ff49d678",
   398 => x"c387f7d8",
   399 => x"496c7cff",
   400 => x"7199ffc3",
   401 => x"f0c3494d",
   402 => x"a9e0c199",
   403 => x"c387cb05",
   404 => x"486c7cff",
   405 => x"66d098c3",
   406 => x"ffc37808",
   407 => x"494a6c7c",
   408 => x"ffc331c8",
   409 => x"714a6c7c",
   410 => x"c84972b2",
   411 => x"7cffc331",
   412 => x"b2714a6c",
   413 => x"31c84972",
   414 => x"6c7cffc3",
   415 => x"ffb2714a",
   416 => x"e0c048d0",
   417 => x"029b7378",
   418 => x"7b7287c2",
   419 => x"4d264875",
   420 => x"4b264c26",
   421 => x"261e4f26",
   422 => x"5b5e0e4f",
   423 => x"86f80e5c",
   424 => x"a6c81e76",
   425 => x"87fdfd49",
   426 => x"4b7086c4",
   427 => x"a8c2486e",
   428 => x"87cac303",
   429 => x"f0c34a73",
   430 => x"aad0c19a",
   431 => x"c187c702",
   432 => x"c205aae0",
   433 => x"497387f8",
   434 => x"c30299c8",
   435 => x"87c6ff87",
   436 => x"9cc34c73",
   437 => x"c105acc2",
   438 => x"66c487cf",
   439 => x"7131c949",
   440 => x"4a66c41e",
   441 => x"c392c8c1",
   442 => x"7249eac9",
   443 => x"ded0fe81",
   444 => x"4966c487",
   445 => x"49e3c01e",
   446 => x"87dbd6ff",
   447 => x"d5ff49d8",
   448 => x"c0c887f0",
   449 => x"daf8c21e",
   450 => x"f3e8fd49",
   451 => x"48d0ff87",
   452 => x"c278e0c0",
   453 => x"d01edaf8",
   454 => x"c8c14a66",
   455 => x"eac9c392",
   456 => x"fe817249",
   457 => x"d087e6cb",
   458 => x"05acc186",
   459 => x"c487cfc1",
   460 => x"31c94966",
   461 => x"66c41e71",
   462 => x"92c8c14a",
   463 => x"49eac9c3",
   464 => x"cffe8172",
   465 => x"f8c287c9",
   466 => x"66c81eda",
   467 => x"92c8c14a",
   468 => x"49eac9c3",
   469 => x"c9fe8172",
   470 => x"66c887f0",
   471 => x"e3c01e49",
   472 => x"f2d4ff49",
   473 => x"ff49d787",
   474 => x"c887c7d4",
   475 => x"f8c21ec0",
   476 => x"e6fd49da",
   477 => x"86d087f4",
   478 => x"c048d0ff",
   479 => x"8ef878e0",
   480 => x"0e87cdfc",
   481 => x"5d5c5b5e",
   482 => x"4d711e0e",
   483 => x"d44cd4ff",
   484 => x"c3487e66",
   485 => x"c506a8b7",
   486 => x"c148c087",
   487 => x"497587e3",
   488 => x"87d2dffe",
   489 => x"66c41e75",
   490 => x"93c8c14b",
   491 => x"83eac9c3",
   492 => x"c3fe4973",
   493 => x"83c887fe",
   494 => x"d0ff4b6b",
   495 => x"78e1c848",
   496 => x"49737cdd",
   497 => x"7199ffc3",
   498 => x"c849737c",
   499 => x"ffc329b7",
   500 => x"737c7199",
   501 => x"29b7d049",
   502 => x"7199ffc3",
   503 => x"d849737c",
   504 => x"7c7129b7",
   505 => x"7c7c7cc0",
   506 => x"7c7c7c7c",
   507 => x"7c7c7c7c",
   508 => x"78e0c07c",
   509 => x"dc1e66c4",
   510 => x"dad2ff49",
   511 => x"7386c887",
   512 => x"c9fa2648",
   513 => x"5b5e0e87",
   514 => x"1e0e5d5c",
   515 => x"d4ff7e71",
   516 => x"c31e6e4b",
   517 => x"fe49facb",
   518 => x"c487d9c2",
   519 => x"9d4d7086",
   520 => x"87c3c302",
   521 => x"bfc2ccc3",
   522 => x"fe496e4c",
   523 => x"ff87c7dd",
   524 => x"c5c848d0",
   525 => x"7bd6c178",
   526 => x"7b154ac0",
   527 => x"e0c082c1",
   528 => x"f504aab7",
   529 => x"48d0ff87",
   530 => x"c5c878c4",
   531 => x"7bd3c178",
   532 => x"78c47bc1",
   533 => x"c1029c74",
   534 => x"f8c287fc",
   535 => x"c0c87eda",
   536 => x"b7c08c4d",
   537 => x"87c603ac",
   538 => x"4da4c0c8",
   539 => x"c5c34cc0",
   540 => x"49bf97cb",
   541 => x"d20299d0",
   542 => x"c31ec087",
   543 => x"fe49facb",
   544 => x"c487c7c5",
   545 => x"4a497086",
   546 => x"c287efc0",
   547 => x"c31edaf8",
   548 => x"fe49facb",
   549 => x"c487f3c4",
   550 => x"4a497086",
   551 => x"c848d0ff",
   552 => x"d4c178c5",
   553 => x"bf976e7b",
   554 => x"c1486e7b",
   555 => x"c17e7080",
   556 => x"f0ff058d",
   557 => x"48d0ff87",
   558 => x"9a7278c4",
   559 => x"c087c505",
   560 => x"87e5c048",
   561 => x"cbc31ec1",
   562 => x"c2fe49fa",
   563 => x"86c487db",
   564 => x"fe059c74",
   565 => x"d0ff87c4",
   566 => x"78c5c848",
   567 => x"c07bd3c1",
   568 => x"c178c47b",
   569 => x"c087c248",
   570 => x"4d262648",
   571 => x"4b264c26",
   572 => x"5e0e4f26",
   573 => x"710e5c5b",
   574 => x"0266cc4b",
   575 => x"c04c87d8",
   576 => x"d8028cf0",
   577 => x"c14a7487",
   578 => x"87d1028a",
   579 => x"87cd028a",
   580 => x"87c9028a",
   581 => x"497387d7",
   582 => x"d087eafb",
   583 => x"c01e7487",
   584 => x"87dff949",
   585 => x"49731e74",
   586 => x"c887d8f9",
   587 => x"87fcfe86",
   588 => x"e5c21e00",
   589 => x"c149bfda",
   590 => x"dee5c2b9",
   591 => x"48d4ff59",
   592 => x"ff78ffc3",
   593 => x"e1c848d0",
   594 => x"48d4ff78",
   595 => x"31c478c1",
   596 => x"d0ff7871",
   597 => x"78e0c048",
   598 => x"00004f26",
   599 => x"ff1e0000",
   600 => x"c487ddc1",
   601 => x"c0c24966",
   602 => x"87cd0299",
   603 => x"c31ee0c3",
   604 => x"ff49f7c8",
   605 => x"c487ecc2",
   606 => x"4966c486",
   607 => x"0299c0c4",
   608 => x"f0c387cd",
   609 => x"f7c8c31e",
   610 => x"d6c2ff49",
   611 => x"c486c487",
   612 => x"ffc14966",
   613 => x"c31e7199",
   614 => x"ff49f7c8",
   615 => x"ff87c4c2",
   616 => x"2687d5c0",
   617 => x"5e0e4f26",
   618 => x"0e5d5c5b",
   619 => x"c086d8ff",
   620 => x"c6cdc37e",
   621 => x"81c249bf",
   622 => x"1e721e71",
   623 => x"dcfd4ac6",
   624 => x"487187f7",
   625 => x"49264a26",
   626 => x"c358a6c8",
   627 => x"49bfc6cd",
   628 => x"1e7181c4",
   629 => x"4ac61e72",
   630 => x"87dddcfd",
   631 => x"4a264871",
   632 => x"a6cc4926",
   633 => x"f7f1c258",
   634 => x"dff049bf",
   635 => x"02987087",
   636 => x"c087f9c9",
   637 => x"c7f049e0",
   638 => x"c2497087",
   639 => x"c059fbf1",
   640 => x"c449744c",
   641 => x"81d0fe91",
   642 => x"49744a69",
   643 => x"bfc6cdc3",
   644 => x"c391c481",
   645 => x"7281d2cd",
   646 => x"d2029a79",
   647 => x"c1497287",
   648 => x"6e9a7189",
   649 => x"7080c148",
   650 => x"059a727e",
   651 => x"c187eeff",
   652 => x"acb7c284",
   653 => x"87c9ff04",
   654 => x"fcc0486e",
   655 => x"c804a8b7",
   656 => x"4cc087ea",
   657 => x"66c44a74",
   658 => x"c392c482",
   659 => x"7482d2cd",
   660 => x"8166c849",
   661 => x"cdc391c4",
   662 => x"4a6a81d2",
   663 => x"b9724969",
   664 => x"cdc34b74",
   665 => x"c483bfc6",
   666 => x"d2cdc393",
   667 => x"72ba6b83",
   668 => x"d4987148",
   669 => x"497458a6",
   670 => x"bfc6cdc3",
   671 => x"c391c481",
   672 => x"6981d2cd",
   673 => x"48a6d47e",
   674 => x"a6d078c0",
   675 => x"4cffc35c",
   676 => x"df4966d0",
   677 => x"e2c60229",
   678 => x"4a66cc87",
   679 => x"d492e0c0",
   680 => x"ffc08266",
   681 => x"70887248",
   682 => x"48a6d84a",
   683 => x"80c478c0",
   684 => x"496e78c0",
   685 => x"e4c029df",
   686 => x"cdc359a6",
   687 => x"78c148c2",
   688 => x"31c34972",
   689 => x"b1722ab7",
   690 => x"c499ffc0",
   691 => x"f3f3c291",
   692 => x"6d85714d",
   693 => x"c0c4494b",
   694 => x"d70299c0",
   695 => x"66e0c087",
   696 => x"87c7c002",
   697 => x"78c080c8",
   698 => x"c387d0c5",
   699 => x"c148cacd",
   700 => x"87c7c578",
   701 => x"0266e0c0",
   702 => x"497387d8",
   703 => x"99c0c0c2",
   704 => x"87c3c002",
   705 => x"6d2bb7d0",
   706 => x"fffffd48",
   707 => x"c07d7098",
   708 => x"cdc387fa",
   709 => x"c002bfca",
   710 => x"487387f2",
   711 => x"c028b7d0",
   712 => x"7058a6e8",
   713 => x"e3c00298",
   714 => x"cecdc387",
   715 => x"e0c049bf",
   716 => x"c00299c0",
   717 => x"497087ca",
   718 => x"99c0e0c0",
   719 => x"87ccc002",
   720 => x"c0c2486d",
   721 => x"7d70b0c0",
   722 => x"4b66e4c0",
   723 => x"c0c84973",
   724 => x"c20299c0",
   725 => x"cdc387c5",
   726 => x"cc4abfce",
   727 => x"c0029ac0",
   728 => x"c0c487cf",
   729 => x"d7c0028a",
   730 => x"c0028a87",
   731 => x"dcc187f8",
   732 => x"74497387",
   733 => x"c291c299",
   734 => x"1181e7f3",
   735 => x"87dbc14b",
   736 => x"99744973",
   737 => x"f3c291c2",
   738 => x"81c181e7",
   739 => x"e0c04b11",
   740 => x"c8c00266",
   741 => x"48a6dc87",
   742 => x"fec078d2",
   743 => x"48a6d887",
   744 => x"c078d2c4",
   745 => x"497387f5",
   746 => x"91c29974",
   747 => x"81e7f3c2",
   748 => x"4b1181c1",
   749 => x"0266e0c0",
   750 => x"dc87c9c0",
   751 => x"d9c148a6",
   752 => x"87d7c078",
   753 => x"c548a6d8",
   754 => x"cec078d9",
   755 => x"74497387",
   756 => x"c291c299",
   757 => x"c181e7f3",
   758 => x"c04b1181",
   759 => x"c00266e0",
   760 => x"497387db",
   761 => x"fcc7b9ff",
   762 => x"487199c0",
   763 => x"bfcecdc3",
   764 => x"d2cdc398",
   765 => x"c49b7458",
   766 => x"d3c0b3c0",
   767 => x"c7497387",
   768 => x"7199c0fc",
   769 => x"cecdc348",
   770 => x"cdc3b0bf",
   771 => x"9b7458d2",
   772 => x"c00266d8",
   773 => x"c31e87ca",
   774 => x"f549c2cd",
   775 => x"86c487c0",
   776 => x"cdc31e73",
   777 => x"f5f449c2",
   778 => x"dc86c487",
   779 => x"cac00266",
   780 => x"cdc31e87",
   781 => x"e5f449c2",
   782 => x"d086c487",
   783 => x"30c14866",
   784 => x"6e58a6d4",
   785 => x"7030c148",
   786 => x"4866d47e",
   787 => x"a6d880c1",
   788 => x"b7e0c058",
   789 => x"f7f804a8",
   790 => x"4c66cc87",
   791 => x"b7c284c1",
   792 => x"dff704ac",
   793 => x"c6cdc387",
   794 => x"7866c448",
   795 => x"268ed8ff",
   796 => x"264c264d",
   797 => x"004f264b",
   798 => x"1e000000",
   799 => x"49724ac0",
   800 => x"cdc391c4",
   801 => x"79ff81d2",
   802 => x"b7c682c1",
   803 => x"87ee04aa",
   804 => x"48c6cdc3",
   805 => x"784040c0",
   806 => x"731e4f26",
   807 => x"f44b711e",
   808 => x"497387c4",
   809 => x"87ecf9fe",
   810 => x"1e87c8ff",
   811 => x"4bc01e73",
   812 => x"49c8f3c2",
   813 => x"7087ceed",
   814 => x"87c40598",
   815 => x"4bd4f3c2",
   816 => x"7387f8fe",
   817 => x"87ebfe48",
   818 => x"4349524f",
   819 => x"20202020",
   820 => x"004d4f52",
   821 => x"204d4f52",
   822 => x"64616f6c",
   823 => x"20676e69",
   824 => x"6c696166",
   825 => x"f4006465",
   826 => x"05f5f2eb",
   827 => x"030c0406",
   828 => x"660a830b",
   829 => x"5a00fc00",
   830 => x"0000da00",
   831 => x"05089480",
   832 => x"02007880",
   833 => x"03000180",
   834 => x"04000980",
   835 => x"01000080",
   836 => x"26089180",
   837 => x"1d000400",
   838 => x"1c000000",
   839 => x"25000000",
   840 => x"1a000c00",
   841 => x"1b000000",
   842 => x"24000000",
   843 => x"12000000",
   844 => x"2e000001",
   845 => x"2d000300",
   846 => x"23000000",
   847 => x"36000000",
   848 => x"21000b00",
   849 => x"2b000000",
   850 => x"2c000000",
   851 => x"22000000",
   852 => x"3d000000",
   853 => x"35006c00",
   854 => x"34000000",
   855 => x"3e000000",
   856 => x"32007500",
   857 => x"33000000",
   858 => x"3c000000",
   859 => x"2a006b00",
   860 => x"46000000",
   861 => x"43000100",
   862 => x"3b007300",
   863 => x"45006900",
   864 => x"3a000900",
   865 => x"42007000",
   866 => x"44007200",
   867 => x"31007400",
   868 => x"55000000",
   869 => x"4d000000",
   870 => x"4b007c00",
   871 => x"7b007a00",
   872 => x"49000000",
   873 => x"4c007100",
   874 => x"54008400",
   875 => x"41007700",
   876 => x"61000000",
   877 => x"5b000000",
   878 => x"52007c00",
   879 => x"f1000000",
   880 => x"59000000",
   881 => x"0e000002",
   882 => x"5d005d00",
   883 => x"4a000000",
   884 => x"16007900",
   885 => x"76000500",
   886 => x"0d000700",
   887 => x"1e000d00",
   888 => x"29000600",
   889 => x"14000000",
   890 => x"15000004",
   891 => x"00000000",
   892 => x"00000040",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
