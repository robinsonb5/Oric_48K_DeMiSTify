library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"eccdc387",
    12 => x"86c0c64e",
    13 => x"49eccdc3",
    14 => x"48f4f7c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087c8e3",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"1e731e4f",
    50 => x"c0029a72",
    51 => x"48c087e7",
    52 => x"a9724bc1",
    53 => x"7287d106",
    54 => x"87c90682",
    55 => x"a9728373",
    56 => x"c387f401",
    57 => x"3ab2c187",
    58 => x"8903a972",
    59 => x"c1078073",
    60 => x"f3052b2a",
    61 => x"264b2687",
    62 => x"1e751e4f",
    63 => x"b7714dc4",
    64 => x"b9ff04a1",
    65 => x"bdc381c1",
    66 => x"a2b77207",
    67 => x"c1baff04",
    68 => x"07bdc182",
    69 => x"c187eefe",
    70 => x"b8ff042d",
    71 => x"2d0780c1",
    72 => x"c1b9ff04",
    73 => x"4d260781",
    74 => x"111e4f26",
    75 => x"08d4ff48",
    76 => x"4866c478",
    77 => x"a6c888c1",
    78 => x"05987058",
    79 => x"4f2687ed",
    80 => x"48d4ff1e",
    81 => x"6878ffc3",
    82 => x"4866c451",
    83 => x"a6c888c1",
    84 => x"05987058",
    85 => x"4f2687eb",
    86 => x"ff1e731e",
    87 => x"ffc34bd4",
    88 => x"c34a6b7b",
    89 => x"496b7bff",
    90 => x"b17232c8",
    91 => x"6b7bffc3",
    92 => x"7131c84a",
    93 => x"7bffc3b2",
    94 => x"32c8496b",
    95 => x"4871b172",
    96 => x"4d2687c4",
    97 => x"4b264c26",
    98 => x"5e0e4f26",
    99 => x"0e5d5c5b",
   100 => x"d4ff4a71",
   101 => x"c349724c",
   102 => x"7c7199ff",
   103 => x"bff4f7c2",
   104 => x"d087c805",
   105 => x"30c94866",
   106 => x"d058a6d4",
   107 => x"29d84966",
   108 => x"7199ffc3",
   109 => x"4966d07c",
   110 => x"ffc329d0",
   111 => x"d07c7199",
   112 => x"29c84966",
   113 => x"7199ffc3",
   114 => x"4966d07c",
   115 => x"7199ffc3",
   116 => x"d049727c",
   117 => x"99ffc329",
   118 => x"4b6c7c71",
   119 => x"4dfff0c9",
   120 => x"05abffc3",
   121 => x"ffc387d0",
   122 => x"c14b6c7c",
   123 => x"87c6028d",
   124 => x"02abffc3",
   125 => x"487387f0",
   126 => x"1e87c7fe",
   127 => x"d4ff49c0",
   128 => x"78ffc348",
   129 => x"c8c381c1",
   130 => x"f104a9b7",
   131 => x"1e4f2687",
   132 => x"87e71e73",
   133 => x"4bdff8c4",
   134 => x"ffc01ec0",
   135 => x"49f7c1f0",
   136 => x"c487e7fd",
   137 => x"05a8c186",
   138 => x"ff87eac0",
   139 => x"ffc348d4",
   140 => x"c0c0c178",
   141 => x"1ec0c0c0",
   142 => x"c1f0e1c0",
   143 => x"c9fd49e9",
   144 => x"7086c487",
   145 => x"87ca0598",
   146 => x"c348d4ff",
   147 => x"48c178ff",
   148 => x"e6fe87cb",
   149 => x"058bc187",
   150 => x"c087fdfe",
   151 => x"87e6fc48",
   152 => x"ff1e731e",
   153 => x"ffc348d4",
   154 => x"c04bd378",
   155 => x"f0ffc01e",
   156 => x"fc49c1c1",
   157 => x"86c487d4",
   158 => x"ca059870",
   159 => x"48d4ff87",
   160 => x"c178ffc3",
   161 => x"fd87cb48",
   162 => x"8bc187f1",
   163 => x"87dbff05",
   164 => x"f1fb48c0",
   165 => x"5b5e0e87",
   166 => x"d4ff0e5c",
   167 => x"87dbfd4c",
   168 => x"c01eeac6",
   169 => x"c8c1f0e1",
   170 => x"87defb49",
   171 => x"a8c186c4",
   172 => x"fe87c802",
   173 => x"48c087ea",
   174 => x"fa87e2c1",
   175 => x"497087da",
   176 => x"99ffffcf",
   177 => x"02a9eac6",
   178 => x"d3fe87c8",
   179 => x"c148c087",
   180 => x"ffc387cb",
   181 => x"4bf1c07c",
   182 => x"7087f4fc",
   183 => x"ebc00298",
   184 => x"c01ec087",
   185 => x"fac1f0ff",
   186 => x"87defa49",
   187 => x"987086c4",
   188 => x"c387d905",
   189 => x"496c7cff",
   190 => x"7c7cffc3",
   191 => x"c0c17c7c",
   192 => x"87c40299",
   193 => x"87d548c1",
   194 => x"87d148c0",
   195 => x"c405abc2",
   196 => x"c848c087",
   197 => x"058bc187",
   198 => x"c087fdfe",
   199 => x"87e4f948",
   200 => x"c21e731e",
   201 => x"c148f4f7",
   202 => x"ff4bc778",
   203 => x"78c248d0",
   204 => x"ff87c8fb",
   205 => x"78c348d0",
   206 => x"e5c01ec0",
   207 => x"49c0c1d0",
   208 => x"c487c7f9",
   209 => x"05a8c186",
   210 => x"c24b87c1",
   211 => x"87c505ab",
   212 => x"f9c048c0",
   213 => x"058bc187",
   214 => x"fc87d0ff",
   215 => x"f7c287f7",
   216 => x"987058f8",
   217 => x"c187cd05",
   218 => x"f0ffc01e",
   219 => x"f849d0c1",
   220 => x"86c487d8",
   221 => x"c348d4ff",
   222 => x"e0c478ff",
   223 => x"fcf7c287",
   224 => x"48d0ff58",
   225 => x"d4ff78c2",
   226 => x"78ffc348",
   227 => x"f5f748c1",
   228 => x"5b5e0e87",
   229 => x"710e5d5c",
   230 => x"4dffc34a",
   231 => x"754cd4ff",
   232 => x"48d0ff7c",
   233 => x"7578c3c4",
   234 => x"c01e727c",
   235 => x"d8c1f0ff",
   236 => x"87d6f749",
   237 => x"987086c4",
   238 => x"c087c502",
   239 => x"87f0c048",
   240 => x"fec37c75",
   241 => x"1ec0c87c",
   242 => x"f54966d4",
   243 => x"86c487dc",
   244 => x"7c757c75",
   245 => x"dad87c75",
   246 => x"7c754be0",
   247 => x"0599496c",
   248 => x"8bc187c5",
   249 => x"7587f305",
   250 => x"48d0ff7c",
   251 => x"48c178c2",
   252 => x"1e87cff6",
   253 => x"ff4ad4ff",
   254 => x"d1c448d0",
   255 => x"7affc378",
   256 => x"f80589c1",
   257 => x"1e4f2687",
   258 => x"4b711e73",
   259 => x"dfcdeec5",
   260 => x"48d4ff4a",
   261 => x"6878ffc3",
   262 => x"a8fec348",
   263 => x"c187c502",
   264 => x"87ed058a",
   265 => x"c5059a72",
   266 => x"c048c087",
   267 => x"9b7387ea",
   268 => x"c887cc02",
   269 => x"49731e66",
   270 => x"c487c5f4",
   271 => x"c887c686",
   272 => x"eefe4966",
   273 => x"48d4ff87",
   274 => x"7878ffc3",
   275 => x"c5059b73",
   276 => x"48d0ff87",
   277 => x"48c178d0",
   278 => x"1e87ebf4",
   279 => x"4a711e73",
   280 => x"d4ff4bc0",
   281 => x"78ffc348",
   282 => x"c448d0ff",
   283 => x"d4ff78c3",
   284 => x"78ffc348",
   285 => x"ffc01e72",
   286 => x"49d1c1f0",
   287 => x"c487cbf4",
   288 => x"05987086",
   289 => x"c0c887cd",
   290 => x"4966cc1e",
   291 => x"c487f8fd",
   292 => x"ff4b7086",
   293 => x"78c248d0",
   294 => x"e9f34873",
   295 => x"5b5e0e87",
   296 => x"c00e5d5c",
   297 => x"f0ffc01e",
   298 => x"f349c9c1",
   299 => x"1ed287dc",
   300 => x"49fcf7c2",
   301 => x"c887d0fd",
   302 => x"c14cc086",
   303 => x"acb7d284",
   304 => x"c287f804",
   305 => x"bf97fcf7",
   306 => x"99c0c349",
   307 => x"05a9c0c1",
   308 => x"c287e7c0",
   309 => x"bf97c3f8",
   310 => x"c231d049",
   311 => x"bf97c4f8",
   312 => x"7232c84a",
   313 => x"c5f8c2b1",
   314 => x"b14abf97",
   315 => x"ffcf4c71",
   316 => x"c19cffff",
   317 => x"c134ca84",
   318 => x"f8c287e7",
   319 => x"49bf97c5",
   320 => x"99c631c1",
   321 => x"97c6f8c2",
   322 => x"b7c74abf",
   323 => x"c2b1722a",
   324 => x"bf97c1f8",
   325 => x"9dcf4d4a",
   326 => x"97c2f8c2",
   327 => x"9ac34abf",
   328 => x"f8c232ca",
   329 => x"4bbf97c3",
   330 => x"b27333c2",
   331 => x"97c4f8c2",
   332 => x"c0c34bbf",
   333 => x"2bb7c69b",
   334 => x"81c2b273",
   335 => x"307148c1",
   336 => x"48c14970",
   337 => x"4d703075",
   338 => x"84c14c72",
   339 => x"c0c89471",
   340 => x"cc06adb7",
   341 => x"b734c187",
   342 => x"b7c0c82d",
   343 => x"f4ff01ad",
   344 => x"f0487487",
   345 => x"5e0e87dc",
   346 => x"0e5d5c5b",
   347 => x"c0c386f8",
   348 => x"78c048e2",
   349 => x"1edaf8c2",
   350 => x"defb49c0",
   351 => x"7086c487",
   352 => x"87c50598",
   353 => x"cec948c0",
   354 => x"c14dc087",
   355 => x"c1fac07e",
   356 => x"f9c249bf",
   357 => x"c8714ad0",
   358 => x"87ceeb4b",
   359 => x"c2059870",
   360 => x"c07ec087",
   361 => x"49bffdf9",
   362 => x"4aecf9c2",
   363 => x"ea4bc871",
   364 => x"987087f8",
   365 => x"c087c205",
   366 => x"c0026e7e",
   367 => x"ffc287fd",
   368 => x"c34dbfe0",
   369 => x"bf9fd8c0",
   370 => x"d6c5487e",
   371 => x"c705a8ea",
   372 => x"e0ffc287",
   373 => x"87ce4dbf",
   374 => x"e9ca486e",
   375 => x"c502a8d5",
   376 => x"c748c087",
   377 => x"f8c287f1",
   378 => x"49751eda",
   379 => x"c487ecf9",
   380 => x"05987086",
   381 => x"48c087c5",
   382 => x"c087dcc7",
   383 => x"49bffdf9",
   384 => x"4aecf9c2",
   385 => x"e94bc871",
   386 => x"987087e0",
   387 => x"c387c805",
   388 => x"c148e2c0",
   389 => x"c087da78",
   390 => x"49bfc1fa",
   391 => x"4ad0f9c2",
   392 => x"e94bc871",
   393 => x"987087c4",
   394 => x"87c5c002",
   395 => x"e6c648c0",
   396 => x"d8c0c387",
   397 => x"c149bf97",
   398 => x"c005a9d5",
   399 => x"c0c387cd",
   400 => x"49bf97d9",
   401 => x"02a9eac2",
   402 => x"c087c5c0",
   403 => x"87c7c648",
   404 => x"97daf8c2",
   405 => x"c3487ebf",
   406 => x"c002a8e9",
   407 => x"486e87ce",
   408 => x"02a8ebc3",
   409 => x"c087c5c0",
   410 => x"87ebc548",
   411 => x"97e5f8c2",
   412 => x"059949bf",
   413 => x"c287ccc0",
   414 => x"bf97e6f8",
   415 => x"02a9c249",
   416 => x"c087c5c0",
   417 => x"87cfc548",
   418 => x"97e7f8c2",
   419 => x"c0c348bf",
   420 => x"4c7058de",
   421 => x"c388c148",
   422 => x"c258e2c0",
   423 => x"bf97e8f8",
   424 => x"c2817549",
   425 => x"bf97e9f8",
   426 => x"7232c84a",
   427 => x"c4c37ea1",
   428 => x"786e48ef",
   429 => x"97eaf8c2",
   430 => x"a6c848bf",
   431 => x"e2c0c358",
   432 => x"d4c202bf",
   433 => x"fdf9c087",
   434 => x"f9c249bf",
   435 => x"c8714aec",
   436 => x"87d6e64b",
   437 => x"c0029870",
   438 => x"48c087c5",
   439 => x"c387f8c3",
   440 => x"4cbfdac0",
   441 => x"5cc3c5c3",
   442 => x"97fff8c2",
   443 => x"31c849bf",
   444 => x"97fef8c2",
   445 => x"49a14abf",
   446 => x"97c0f9c2",
   447 => x"32d04abf",
   448 => x"c249a172",
   449 => x"bf97c1f9",
   450 => x"7232d84a",
   451 => x"66c449a1",
   452 => x"efc4c391",
   453 => x"c4c381bf",
   454 => x"f9c259f7",
   455 => x"4abf97c7",
   456 => x"f9c232c8",
   457 => x"4bbf97c6",
   458 => x"f9c24aa2",
   459 => x"4bbf97c8",
   460 => x"a27333d0",
   461 => x"c9f9c24a",
   462 => x"cf4bbf97",
   463 => x"7333d89b",
   464 => x"c4c34aa2",
   465 => x"c4c35afb",
   466 => x"c24abff7",
   467 => x"c392748a",
   468 => x"7248fbc4",
   469 => x"cac178a1",
   470 => x"ecf8c287",
   471 => x"c849bf97",
   472 => x"ebf8c231",
   473 => x"a14abf97",
   474 => x"eac0c349",
   475 => x"e6c0c359",
   476 => x"31c549bf",
   477 => x"c981ffc7",
   478 => x"c3c5c329",
   479 => x"f1f8c259",
   480 => x"c84abf97",
   481 => x"f0f8c232",
   482 => x"a24bbf97",
   483 => x"9266c44a",
   484 => x"c4c3826e",
   485 => x"c4c35aff",
   486 => x"78c048f7",
   487 => x"48f3c4c3",
   488 => x"c378a172",
   489 => x"c348c3c5",
   490 => x"78bff7c4",
   491 => x"48c7c5c3",
   492 => x"bffbc4c3",
   493 => x"e2c0c378",
   494 => x"c9c002bf",
   495 => x"c4487487",
   496 => x"c07e7030",
   497 => x"c4c387c9",
   498 => x"c448bfff",
   499 => x"c37e7030",
   500 => x"6e48e6c0",
   501 => x"f848c178",
   502 => x"264d268e",
   503 => x"264b264c",
   504 => x"5b5e0e4f",
   505 => x"710e5d5c",
   506 => x"e2c0c34a",
   507 => x"87cb02bf",
   508 => x"2bc74b72",
   509 => x"ffc14c72",
   510 => x"7287c99c",
   511 => x"722bc84b",
   512 => x"9cffc34c",
   513 => x"bfefc4c3",
   514 => x"f9f9c083",
   515 => x"d902abbf",
   516 => x"fdf9c087",
   517 => x"daf8c25b",
   518 => x"f049731e",
   519 => x"86c487fd",
   520 => x"c5059870",
   521 => x"c048c087",
   522 => x"c0c387e6",
   523 => x"d202bfe2",
   524 => x"c4497487",
   525 => x"daf8c291",
   526 => x"cf4d6981",
   527 => x"ffffffff",
   528 => x"7487cb9d",
   529 => x"c291c249",
   530 => x"9f81daf8",
   531 => x"48754d69",
   532 => x"0e87c6fe",
   533 => x"5d5c5b5e",
   534 => x"4d711e0e",
   535 => x"49c11ec0",
   536 => x"c487fed0",
   537 => x"9c4c7086",
   538 => x"87c2c102",
   539 => x"4aeac0c3",
   540 => x"dfff4975",
   541 => x"987087d9",
   542 => x"87f2c002",
   543 => x"49754a74",
   544 => x"dfff4bcb",
   545 => x"987087fe",
   546 => x"87e2c002",
   547 => x"9c741ec0",
   548 => x"c487c702",
   549 => x"78c048a6",
   550 => x"a6c487c5",
   551 => x"c478c148",
   552 => x"fccf4966",
   553 => x"7086c487",
   554 => x"fe059c4c",
   555 => x"487487fe",
   556 => x"87e5fc26",
   557 => x"5c5b5e0e",
   558 => x"86f80e5d",
   559 => x"059b4b71",
   560 => x"48c087c5",
   561 => x"c887ddc2",
   562 => x"7dc04da3",
   563 => x"c70266d8",
   564 => x"9766d887",
   565 => x"87c505bf",
   566 => x"c7c248c0",
   567 => x"4966d887",
   568 => x"7087f0fd",
   569 => x"c1026e7e",
   570 => x"496e87f8",
   571 => x"7d6981dc",
   572 => x"81da496e",
   573 => x"9f4ca3c4",
   574 => x"c0c37c69",
   575 => x"d002bfe2",
   576 => x"d4496e87",
   577 => x"49699f81",
   578 => x"ffffc04a",
   579 => x"c232d09a",
   580 => x"724ac087",
   581 => x"806c4849",
   582 => x"7bc07c70",
   583 => x"6c49a3cc",
   584 => x"49a3d079",
   585 => x"a6c479c0",
   586 => x"d478c048",
   587 => x"66c44aa3",
   588 => x"7291c849",
   589 => x"41c049a1",
   590 => x"66c4796c",
   591 => x"c880c148",
   592 => x"b7c658a6",
   593 => x"e2ff04a8",
   594 => x"c94a6d87",
   595 => x"c049722a",
   596 => x"ddff4af0",
   597 => x"4a7087ef",
   598 => x"49a3c4c1",
   599 => x"486e7972",
   600 => x"48c087c2",
   601 => x"f0f98ef8",
   602 => x"5b5e0e87",
   603 => x"710e5d5c",
   604 => x"f9f9c04c",
   605 => x"7478ff48",
   606 => x"cac1029c",
   607 => x"49a4c887",
   608 => x"c2c10269",
   609 => x"4a66d087",
   610 => x"d482496c",
   611 => x"66d05aa6",
   612 => x"c0c3b94d",
   613 => x"ff4abfde",
   614 => x"719972ba",
   615 => x"e4c00299",
   616 => x"4ba4c487",
   617 => x"f8f8496b",
   618 => x"c37b7087",
   619 => x"49bfdac0",
   620 => x"7c71816c",
   621 => x"c0c3b975",
   622 => x"ff4abfde",
   623 => x"719972ba",
   624 => x"dcff0599",
   625 => x"f87c7587",
   626 => x"731e87cf",
   627 => x"9b4b711e",
   628 => x"c887c702",
   629 => x"056949a3",
   630 => x"48c087c5",
   631 => x"c387ebc0",
   632 => x"4abff3c4",
   633 => x"6949a3c4",
   634 => x"c389c249",
   635 => x"91bfdac0",
   636 => x"c34aa271",
   637 => x"49bfdec0",
   638 => x"a271996b",
   639 => x"1e66c84a",
   640 => x"d6e94972",
   641 => x"7086c487",
   642 => x"d0f74849",
   643 => x"1e731e87",
   644 => x"029b4b71",
   645 => x"a3c887c7",
   646 => x"c5056949",
   647 => x"c048c087",
   648 => x"c4c387eb",
   649 => x"c44abff3",
   650 => x"496949a3",
   651 => x"c0c389c2",
   652 => x"7191bfda",
   653 => x"c0c34aa2",
   654 => x"6b49bfde",
   655 => x"4aa27199",
   656 => x"721e66c8",
   657 => x"87c9e549",
   658 => x"497086c4",
   659 => x"87cdf648",
   660 => x"5c5b5e0e",
   661 => x"86f80e5d",
   662 => x"a6c44b71",
   663 => x"c878ff48",
   664 => x"4d6949a3",
   665 => x"a3d44cc0",
   666 => x"c849744a",
   667 => x"49a17291",
   668 => x"66d84969",
   669 => x"70887148",
   670 => x"a966d87e",
   671 => x"6e87ca01",
   672 => x"87c506ad",
   673 => x"6e5ca6c8",
   674 => x"c684c14d",
   675 => x"ff04acb7",
   676 => x"66c487d4",
   677 => x"f48ef848",
   678 => x"5e0e87ff",
   679 => x"0e5d5c5b",
   680 => x"a6c886ec",
   681 => x"48a6c859",
   682 => x"ffffffc1",
   683 => x"c478ffff",
   684 => x"c078ff80",
   685 => x"c44cc04d",
   686 => x"83d44b66",
   687 => x"91c84974",
   688 => x"7549a173",
   689 => x"7392c84a",
   690 => x"49697ea2",
   691 => x"d489bf6e",
   692 => x"ad7459a6",
   693 => x"d087c605",
   694 => x"bf6e48a6",
   695 => x"4866d078",
   696 => x"04a8b7c0",
   697 => x"66d087cf",
   698 => x"a966c849",
   699 => x"d087c603",
   700 => x"a6cc5ca6",
   701 => x"c684c159",
   702 => x"fe04acb7",
   703 => x"85c187f9",
   704 => x"04adb7c6",
   705 => x"cc87eefe",
   706 => x"8eec4866",
   707 => x"0e87caf3",
   708 => x"5d5c5b5e",
   709 => x"7186f00e",
   710 => x"66e0c04b",
   711 => x"732cc94c",
   712 => x"e1c3029b",
   713 => x"49a3c887",
   714 => x"d9c30269",
   715 => x"49a3d087",
   716 => x"7966e0c0",
   717 => x"02ac7e6b",
   718 => x"c387cbc3",
   719 => x"49bfdec0",
   720 => x"4a71b9ff",
   721 => x"48719a74",
   722 => x"a6cc986e",
   723 => x"4da3c458",
   724 => x"6d48a6c4",
   725 => x"aa66c878",
   726 => x"7487c505",
   727 => x"87d1c27b",
   728 => x"49731e72",
   729 => x"c487e9fb",
   730 => x"487e7086",
   731 => x"04a8b7c0",
   732 => x"a3d487d0",
   733 => x"c8496e4a",
   734 => x"49a17291",
   735 => x"7d697b21",
   736 => x"7bc087c7",
   737 => x"6949a3cc",
   738 => x"1e66c87d",
   739 => x"fffa4973",
   740 => x"7086c487",
   741 => x"a3c4c17e",
   742 => x"48a6cc49",
   743 => x"66c87869",
   744 => x"a866cc48",
   745 => x"6e87c906",
   746 => x"a8b7c048",
   747 => x"87e0c004",
   748 => x"b7c0486e",
   749 => x"ecc004a8",
   750 => x"4aa3d487",
   751 => x"91c8496e",
   752 => x"c849a172",
   753 => x"88694866",
   754 => x"66cc4970",
   755 => x"87d506a9",
   756 => x"c5fb4973",
   757 => x"d4497087",
   758 => x"91c84aa3",
   759 => x"c849a172",
   760 => x"66c44166",
   761 => x"748c6b79",
   762 => x"49731e49",
   763 => x"c487faf5",
   764 => x"66e0c086",
   765 => x"99ffc749",
   766 => x"c287cb02",
   767 => x"731edaf8",
   768 => x"87c6f749",
   769 => x"8ef086c4",
   770 => x"1e87ceef",
   771 => x"4b711e73",
   772 => x"e4c0029b",
   773 => x"c7c5c387",
   774 => x"c24a735b",
   775 => x"dac0c38a",
   776 => x"c39249bf",
   777 => x"48bff3c4",
   778 => x"c5c38072",
   779 => x"487158cb",
   780 => x"c0c330c4",
   781 => x"edc058ea",
   782 => x"c3c5c387",
   783 => x"f7c4c348",
   784 => x"c5c378bf",
   785 => x"c4c348c7",
   786 => x"c378bffb",
   787 => x"02bfe2c0",
   788 => x"c0c387c9",
   789 => x"c449bfda",
   790 => x"c387c731",
   791 => x"49bfffc4",
   792 => x"c0c331c4",
   793 => x"f4ed59ea",
   794 => x"5b5e0e87",
   795 => x"4a710e5c",
   796 => x"9a724bc0",
   797 => x"87e1c002",
   798 => x"9f49a2da",
   799 => x"c0c34b69",
   800 => x"cf02bfe2",
   801 => x"49a2d487",
   802 => x"4c49699f",
   803 => x"9cffffc0",
   804 => x"87c234d0",
   805 => x"49744cc0",
   806 => x"fd4973b3",
   807 => x"faec87ed",
   808 => x"5b5e0e87",
   809 => x"f40e5d5c",
   810 => x"c04a7186",
   811 => x"029a727e",
   812 => x"f8c287d8",
   813 => x"78c048d6",
   814 => x"48cef8c2",
   815 => x"bfc7c5c3",
   816 => x"d2f8c278",
   817 => x"c3c5c348",
   818 => x"c0c378bf",
   819 => x"50c048f7",
   820 => x"bfe6c0c3",
   821 => x"d6f8c249",
   822 => x"aa714abf",
   823 => x"87c0c403",
   824 => x"99cf4972",
   825 => x"87e1c005",
   826 => x"1edaf8c2",
   827 => x"bfcef8c2",
   828 => x"cef8c249",
   829 => x"78a1c148",
   830 => x"deddff71",
   831 => x"c086c487",
   832 => x"c248f5f9",
   833 => x"cc78daf8",
   834 => x"f5f9c087",
   835 => x"e0c048bf",
   836 => x"f9f9c080",
   837 => x"d6f8c258",
   838 => x"80c148bf",
   839 => x"58daf8c2",
   840 => x"000e7527",
   841 => x"bf97bf00",
   842 => x"c2029d4d",
   843 => x"e5c387e2",
   844 => x"dbc202ad",
   845 => x"f5f9c087",
   846 => x"a3cb4bbf",
   847 => x"cf4c1149",
   848 => x"d2c105ac",
   849 => x"df497587",
   850 => x"cd89c199",
   851 => x"eac0c391",
   852 => x"4aa3c181",
   853 => x"a3c35112",
   854 => x"c551124a",
   855 => x"51124aa3",
   856 => x"124aa3c7",
   857 => x"4aa3c951",
   858 => x"a3ce5112",
   859 => x"d051124a",
   860 => x"51124aa3",
   861 => x"124aa3d2",
   862 => x"4aa3d451",
   863 => x"a3d65112",
   864 => x"d851124a",
   865 => x"51124aa3",
   866 => x"124aa3dc",
   867 => x"4aa3de51",
   868 => x"7ec15112",
   869 => x"7487f9c0",
   870 => x"0599c849",
   871 => x"7487eac0",
   872 => x"0599d049",
   873 => x"66dc87d0",
   874 => x"87cac002",
   875 => x"66dc4973",
   876 => x"0298700f",
   877 => x"056e87d3",
   878 => x"c387c6c0",
   879 => x"c048eac0",
   880 => x"f5f9c050",
   881 => x"e7c248bf",
   882 => x"f7c0c387",
   883 => x"7e50c048",
   884 => x"bfe6c0c3",
   885 => x"d6f8c249",
   886 => x"aa714abf",
   887 => x"87c0fc04",
   888 => x"bfc7c5c3",
   889 => x"87c8c005",
   890 => x"bfe2c0c3",
   891 => x"87fec102",
   892 => x"48f9f9c0",
   893 => x"f8c278ff",
   894 => x"e749bfd2",
   895 => x"497087e3",
   896 => x"59d6f8c2",
   897 => x"c248a6c4",
   898 => x"78bfd2f8",
   899 => x"bfe2c0c3",
   900 => x"87d8c002",
   901 => x"cf4966c4",
   902 => x"f8ffffff",
   903 => x"c002a999",
   904 => x"4dc087c5",
   905 => x"c187e1c0",
   906 => x"87dcc04d",
   907 => x"cf4966c4",
   908 => x"a999f8ff",
   909 => x"87c8c002",
   910 => x"c048a6c8",
   911 => x"87c5c078",
   912 => x"c148a6c8",
   913 => x"4d66c878",
   914 => x"c0059d75",
   915 => x"66c487e0",
   916 => x"c389c249",
   917 => x"4abfdac0",
   918 => x"f3c4c391",
   919 => x"f8c24abf",
   920 => x"a17248ce",
   921 => x"d6f8c278",
   922 => x"f978c048",
   923 => x"48c087e2",
   924 => x"e4e58ef4",
   925 => x"00000087",
   926 => x"ffffff00",
   927 => x"000e85ff",
   928 => x"000e8e00",
   929 => x"54414600",
   930 => x"20203233",
   931 => x"41460020",
   932 => x"20363154",
   933 => x"1e002020",
   934 => x"c348d4ff",
   935 => x"486878ff",
   936 => x"ff1e4f26",
   937 => x"ffc348d4",
   938 => x"48d0ff78",
   939 => x"ff78e1c8",
   940 => x"78d448d4",
   941 => x"48cbc5c3",
   942 => x"50bfd4ff",
   943 => x"ff1e4f26",
   944 => x"e0c048d0",
   945 => x"1e4f2678",
   946 => x"7087ccff",
   947 => x"c6029949",
   948 => x"a9fbc087",
   949 => x"7187f105",
   950 => x"0e4f2648",
   951 => x"0e5c5b5e",
   952 => x"4cc04b71",
   953 => x"7087f0fe",
   954 => x"c0029949",
   955 => x"ecc087f9",
   956 => x"f2c002a9",
   957 => x"a9fbc087",
   958 => x"87ebc002",
   959 => x"acb766cc",
   960 => x"d087c703",
   961 => x"87c20266",
   962 => x"99715371",
   963 => x"c187c202",
   964 => x"87c3fe84",
   965 => x"02994970",
   966 => x"ecc087cd",
   967 => x"87c702a9",
   968 => x"05a9fbc0",
   969 => x"d087d5ff",
   970 => x"87c30266",
   971 => x"c07b97c0",
   972 => x"c405a9ec",
   973 => x"c54a7487",
   974 => x"c04a7487",
   975 => x"48728a0a",
   976 => x"4d2687c2",
   977 => x"4b264c26",
   978 => x"fd1e4f26",
   979 => x"497087c9",
   980 => x"a9b7f0c0",
   981 => x"c087ca04",
   982 => x"01a9b7f9",
   983 => x"f0c087c3",
   984 => x"b7c1c189",
   985 => x"87ca04a9",
   986 => x"a9b7dac1",
   987 => x"c087c301",
   988 => x"487189f7",
   989 => x"5e0e4f26",
   990 => x"710e5c5b",
   991 => x"4cd4ff4a",
   992 => x"eac04972",
   993 => x"9b4b7087",
   994 => x"c187c202",
   995 => x"48d0ff8b",
   996 => x"c178c5c8",
   997 => x"49737cd5",
   998 => x"e4c231c6",
   999 => x"4abf97f0",
  1000 => x"70b07148",
  1001 => x"48d0ff7c",
  1002 => x"487378c4",
  1003 => x"0e87d5fe",
  1004 => x"5d5c5b5e",
  1005 => x"7186f80e",
  1006 => x"fb7ec04c",
  1007 => x"4bc087e4",
  1008 => x"97dcc1c1",
  1009 => x"a9c049bf",
  1010 => x"fb87cf04",
  1011 => x"83c187f9",
  1012 => x"97dcc1c1",
  1013 => x"06ab49bf",
  1014 => x"c1c187f1",
  1015 => x"02bf97dc",
  1016 => x"f2fa87cf",
  1017 => x"99497087",
  1018 => x"c087c602",
  1019 => x"f105a9ec",
  1020 => x"fa4bc087",
  1021 => x"4d7087e1",
  1022 => x"c887dcfa",
  1023 => x"d6fa58a6",
  1024 => x"c14a7087",
  1025 => x"49a4c883",
  1026 => x"ad496997",
  1027 => x"c087c702",
  1028 => x"c005adff",
  1029 => x"a4c987e7",
  1030 => x"49699749",
  1031 => x"02a966c4",
  1032 => x"c04887c7",
  1033 => x"d405a8ff",
  1034 => x"49a4ca87",
  1035 => x"aa496997",
  1036 => x"c087c602",
  1037 => x"c405aaff",
  1038 => x"d07ec187",
  1039 => x"adecc087",
  1040 => x"c087c602",
  1041 => x"c405adfb",
  1042 => x"c14bc087",
  1043 => x"fe026e7e",
  1044 => x"e9f987e1",
  1045 => x"f8487387",
  1046 => x"87e6fb8e",
  1047 => x"5b5e0e00",
  1048 => x"1e0e5d5c",
  1049 => x"4cc04b71",
  1050 => x"c004ab4d",
  1051 => x"fec087e8",
  1052 => x"9d751eef",
  1053 => x"c087c402",
  1054 => x"c187c24a",
  1055 => x"f049724a",
  1056 => x"86c487df",
  1057 => x"84c17e70",
  1058 => x"87c2056e",
  1059 => x"85c14c73",
  1060 => x"ff06ac73",
  1061 => x"486e87d8",
  1062 => x"264d2626",
  1063 => x"264b264c",
  1064 => x"5b5e0e4f",
  1065 => x"1e0e5d5c",
  1066 => x"de494c71",
  1067 => x"e5c5c391",
  1068 => x"9785714d",
  1069 => x"ddc1026d",
  1070 => x"d0c5c387",
  1071 => x"82744abf",
  1072 => x"d8fe4972",
  1073 => x"6e7e7087",
  1074 => x"87f3c002",
  1075 => x"4bd8c5c3",
  1076 => x"49cb4a6e",
  1077 => x"87d0fffe",
  1078 => x"93cb4b74",
  1079 => x"83f7e4c1",
  1080 => x"c4c183c4",
  1081 => x"49747bda",
  1082 => x"87d9c2c1",
  1083 => x"c5c37b75",
  1084 => x"49bf97e4",
  1085 => x"d8c5c31e",
  1086 => x"f5dfc149",
  1087 => x"7486c487",
  1088 => x"c0c2c149",
  1089 => x"c149c087",
  1090 => x"c387dfc3",
  1091 => x"c048ccc5",
  1092 => x"dd49c178",
  1093 => x"fd2687cb",
  1094 => x"6f4c87ff",
  1095 => x"6e696461",
  1096 => x"2e2e2e67",
  1097 => x"5b5e0e00",
  1098 => x"4b710e5c",
  1099 => x"d0c5c34a",
  1100 => x"497282bf",
  1101 => x"7087e6fc",
  1102 => x"c4029c4c",
  1103 => x"e8ec4987",
  1104 => x"d0c5c387",
  1105 => x"c178c048",
  1106 => x"87d5dc49",
  1107 => x"0e87ccfd",
  1108 => x"5d5c5b5e",
  1109 => x"c286f40e",
  1110 => x"c04ddaf8",
  1111 => x"48a6c44c",
  1112 => x"c5c378c0",
  1113 => x"c049bfd0",
  1114 => x"c1c106a9",
  1115 => x"daf8c287",
  1116 => x"c0029848",
  1117 => x"fec087f8",
  1118 => x"66c81eef",
  1119 => x"c487c702",
  1120 => x"78c048a6",
  1121 => x"a6c487c5",
  1122 => x"c478c148",
  1123 => x"d0ec4966",
  1124 => x"7086c487",
  1125 => x"c484c14d",
  1126 => x"80c14866",
  1127 => x"c358a6c8",
  1128 => x"49bfd0c5",
  1129 => x"87c603ac",
  1130 => x"ff059d75",
  1131 => x"4cc087c8",
  1132 => x"c3029d75",
  1133 => x"fec087e0",
  1134 => x"66c81eef",
  1135 => x"cc87c702",
  1136 => x"78c048a6",
  1137 => x"a6cc87c5",
  1138 => x"cc78c148",
  1139 => x"d0eb4966",
  1140 => x"7086c487",
  1141 => x"c2026e7e",
  1142 => x"496e87e9",
  1143 => x"699781cb",
  1144 => x"0299d049",
  1145 => x"c187d6c1",
  1146 => x"744ae5c4",
  1147 => x"c191cb49",
  1148 => x"7281f7e4",
  1149 => x"c381c879",
  1150 => x"497451ff",
  1151 => x"c5c391de",
  1152 => x"85714de5",
  1153 => x"7d97c1c2",
  1154 => x"c049a5c1",
  1155 => x"c0c351e0",
  1156 => x"02bf97ea",
  1157 => x"84c187d2",
  1158 => x"c34ba5c2",
  1159 => x"db4aeac0",
  1160 => x"c3fafe49",
  1161 => x"87dbc187",
  1162 => x"c049a5cd",
  1163 => x"c284c151",
  1164 => x"4a6e4ba5",
  1165 => x"f9fe49cb",
  1166 => x"c6c187ee",
  1167 => x"e1c2c187",
  1168 => x"cb49744a",
  1169 => x"f7e4c191",
  1170 => x"c3797281",
  1171 => x"bf97eac0",
  1172 => x"7487d802",
  1173 => x"c191de49",
  1174 => x"e5c5c384",
  1175 => x"c383714b",
  1176 => x"dd4aeac0",
  1177 => x"fff8fe49",
  1178 => x"7487d887",
  1179 => x"c393de4b",
  1180 => x"cb83e5c5",
  1181 => x"51c049a3",
  1182 => x"6e7384c1",
  1183 => x"fe49cb4a",
  1184 => x"c487e5f8",
  1185 => x"80c14866",
  1186 => x"c758a6c8",
  1187 => x"c5c003ac",
  1188 => x"fc056e87",
  1189 => x"487487e0",
  1190 => x"fcf78ef4",
  1191 => x"1e731e87",
  1192 => x"cb494b71",
  1193 => x"f7e4c191",
  1194 => x"4aa1c881",
  1195 => x"48f0e4c2",
  1196 => x"a1c95012",
  1197 => x"dcc1c14a",
  1198 => x"ca501248",
  1199 => x"e4c5c381",
  1200 => x"c3501148",
  1201 => x"bf97e4c5",
  1202 => x"49c01e49",
  1203 => x"87e2d8c1",
  1204 => x"48ccc5c3",
  1205 => x"49c178de",
  1206 => x"2687c6d6",
  1207 => x"1e87fef6",
  1208 => x"cb494a71",
  1209 => x"f7e4c191",
  1210 => x"1181c881",
  1211 => x"d0c5c348",
  1212 => x"d0c5c358",
  1213 => x"c178c048",
  1214 => x"87e5d549",
  1215 => x"c01e4f26",
  1216 => x"e5fbc049",
  1217 => x"1e4f2687",
  1218 => x"d2029971",
  1219 => x"cce6c187",
  1220 => x"f750c048",
  1221 => x"dfcbc180",
  1222 => x"f0e4c140",
  1223 => x"c187ce78",
  1224 => x"c148c8e6",
  1225 => x"fc78e9e4",
  1226 => x"fecbc180",
  1227 => x"0e4f2678",
  1228 => x"0e5c5b5e",
  1229 => x"cb4a4c71",
  1230 => x"f7e4c192",
  1231 => x"49a2c882",
  1232 => x"974ba2c9",
  1233 => x"971e4b6b",
  1234 => x"ca1e4969",
  1235 => x"c0491282",
  1236 => x"c087e0e6",
  1237 => x"87c9d449",
  1238 => x"f8c04974",
  1239 => x"8ef887e7",
  1240 => x"1e87f8f4",
  1241 => x"4b711e73",
  1242 => x"87c3ff49",
  1243 => x"fefe4973",
  1244 => x"87e9f487",
  1245 => x"711e731e",
  1246 => x"4aa3c64b",
  1247 => x"c187db02",
  1248 => x"87d6028a",
  1249 => x"dac1028a",
  1250 => x"c0028a87",
  1251 => x"028a87fc",
  1252 => x"8a87e1c0",
  1253 => x"c187cb02",
  1254 => x"49c787db",
  1255 => x"c187c0fd",
  1256 => x"c5c387de",
  1257 => x"c102bfd0",
  1258 => x"c14887cb",
  1259 => x"d4c5c388",
  1260 => x"87c1c158",
  1261 => x"bfd4c5c3",
  1262 => x"87f9c002",
  1263 => x"bfd0c5c3",
  1264 => x"c380c148",
  1265 => x"c058d4c5",
  1266 => x"c5c387eb",
  1267 => x"c649bfd0",
  1268 => x"d4c5c389",
  1269 => x"a9b7c059",
  1270 => x"c387da03",
  1271 => x"c048d0c5",
  1272 => x"c387d278",
  1273 => x"02bfd4c5",
  1274 => x"c5c387cb",
  1275 => x"c648bfd0",
  1276 => x"d4c5c380",
  1277 => x"d149c058",
  1278 => x"497387e7",
  1279 => x"87c5f6c0",
  1280 => x"0e87daf2",
  1281 => x"0e5c5b5e",
  1282 => x"66cc4c71",
  1283 => x"cb4b741e",
  1284 => x"f7e4c193",
  1285 => x"4aa3c483",
  1286 => x"f2fe496a",
  1287 => x"cac187da",
  1288 => x"a3c87bdd",
  1289 => x"5166d449",
  1290 => x"d849a3c9",
  1291 => x"a3ca5166",
  1292 => x"5166dc49",
  1293 => x"87e3f126",
  1294 => x"5c5b5e0e",
  1295 => x"d0ff0e5d",
  1296 => x"59a6d886",
  1297 => x"c048a6c4",
  1298 => x"c180c478",
  1299 => x"c47866c4",
  1300 => x"c478c180",
  1301 => x"c378c180",
  1302 => x"c148d4c5",
  1303 => x"ccc5c378",
  1304 => x"a8de48bf",
  1305 => x"f387cb05",
  1306 => x"497087e5",
  1307 => x"ce59a6c8",
  1308 => x"ede887f8",
  1309 => x"87cfe987",
  1310 => x"7087dce8",
  1311 => x"acfbc04c",
  1312 => x"87d0c102",
  1313 => x"c10566d4",
  1314 => x"1ec087c2",
  1315 => x"c11ec11e",
  1316 => x"c01edae6",
  1317 => x"87ebfd49",
  1318 => x"4a66d0c1",
  1319 => x"496a82c4",
  1320 => x"517481c7",
  1321 => x"1ed81ec1",
  1322 => x"81c8496a",
  1323 => x"d887ece8",
  1324 => x"66c4c186",
  1325 => x"01a8c048",
  1326 => x"a6c487c7",
  1327 => x"ce78c148",
  1328 => x"66c4c187",
  1329 => x"cc88c148",
  1330 => x"87c358a6",
  1331 => x"cc87f8e7",
  1332 => x"78c248a6",
  1333 => x"cd029c74",
  1334 => x"66c487cc",
  1335 => x"66c8c148",
  1336 => x"c1cd03a8",
  1337 => x"48a6d887",
  1338 => x"eae678c0",
  1339 => x"c14c7087",
  1340 => x"c205acd0",
  1341 => x"66d887d6",
  1342 => x"87cee97e",
  1343 => x"a6dc4970",
  1344 => x"87d3e659",
  1345 => x"ecc04c70",
  1346 => x"eac105ac",
  1347 => x"4966c487",
  1348 => x"c0c191cb",
  1349 => x"a1c48166",
  1350 => x"c84d6a4a",
  1351 => x"66d84aa1",
  1352 => x"dfcbc152",
  1353 => x"87efe579",
  1354 => x"029c4c70",
  1355 => x"fbc087d8",
  1356 => x"87d202ac",
  1357 => x"dee55574",
  1358 => x"9c4c7087",
  1359 => x"c087c702",
  1360 => x"ff05acfb",
  1361 => x"e0c087ee",
  1362 => x"55c1c255",
  1363 => x"d47d97c0",
  1364 => x"a96e4966",
  1365 => x"c487db05",
  1366 => x"66c84866",
  1367 => x"87ca04a8",
  1368 => x"c14866c4",
  1369 => x"58a6c880",
  1370 => x"66c887c8",
  1371 => x"cc88c148",
  1372 => x"e2e458a6",
  1373 => x"c14c7087",
  1374 => x"c805acd0",
  1375 => x"4866d087",
  1376 => x"a6d480c1",
  1377 => x"acd0c158",
  1378 => x"87eafd02",
  1379 => x"d448a6dc",
  1380 => x"66d87866",
  1381 => x"a866dc48",
  1382 => x"87dcc905",
  1383 => x"48a6e0c0",
  1384 => x"c478f0c0",
  1385 => x"7866cc80",
  1386 => x"78c080c4",
  1387 => x"c048747e",
  1388 => x"f0c088fb",
  1389 => x"987058a6",
  1390 => x"87d7c802",
  1391 => x"c088cb48",
  1392 => x"7058a6f0",
  1393 => x"e9c00298",
  1394 => x"88c94887",
  1395 => x"58a6f0c0",
  1396 => x"c3029870",
  1397 => x"c44887e1",
  1398 => x"a6f0c088",
  1399 => x"02987058",
  1400 => x"c14887d6",
  1401 => x"a6f0c088",
  1402 => x"02987058",
  1403 => x"c787c8c3",
  1404 => x"e0c087db",
  1405 => x"78c048a6",
  1406 => x"c14866cc",
  1407 => x"58a6d080",
  1408 => x"7087d4e2",
  1409 => x"acecc04c",
  1410 => x"c087d502",
  1411 => x"c60266e0",
  1412 => x"a6e4c087",
  1413 => x"7487c95c",
  1414 => x"88f0c048",
  1415 => x"58a6e8c0",
  1416 => x"02acecc0",
  1417 => x"eee187cc",
  1418 => x"c04c7087",
  1419 => x"ff05acec",
  1420 => x"e0c087f4",
  1421 => x"66d41e66",
  1422 => x"ecc01e49",
  1423 => x"e6c11e66",
  1424 => x"66d41eda",
  1425 => x"87fbf649",
  1426 => x"1eca1ec0",
  1427 => x"cb4966dc",
  1428 => x"66d8c191",
  1429 => x"48a6d881",
  1430 => x"d878a1c4",
  1431 => x"e149bf66",
  1432 => x"86d887f9",
  1433 => x"06a8b7c0",
  1434 => x"c187c7c1",
  1435 => x"c81ede1e",
  1436 => x"e149bf66",
  1437 => x"86c887e5",
  1438 => x"c0484970",
  1439 => x"e4c08808",
  1440 => x"b7c058a6",
  1441 => x"e9c006a8",
  1442 => x"66e0c087",
  1443 => x"a8b7dd48",
  1444 => x"6e87df03",
  1445 => x"e0c049bf",
  1446 => x"e0c08166",
  1447 => x"c1496651",
  1448 => x"81bf6e81",
  1449 => x"c051c1c2",
  1450 => x"c24966e0",
  1451 => x"81bf6e81",
  1452 => x"7ec151c0",
  1453 => x"e287dcc4",
  1454 => x"e4c087d0",
  1455 => x"c9e258a6",
  1456 => x"a6e8c087",
  1457 => x"a8ecc058",
  1458 => x"87cbc005",
  1459 => x"48a6e4c0",
  1460 => x"7866e0c0",
  1461 => x"ff87c4c0",
  1462 => x"c487fcde",
  1463 => x"91cb4966",
  1464 => x"4866c0c1",
  1465 => x"7e708071",
  1466 => x"82c84a6e",
  1467 => x"81ca496e",
  1468 => x"5166e0c0",
  1469 => x"4966e4c0",
  1470 => x"e0c081c1",
  1471 => x"48c18966",
  1472 => x"49703071",
  1473 => x"977189c1",
  1474 => x"c1c9c37a",
  1475 => x"e0c049bf",
  1476 => x"6a972966",
  1477 => x"9871484a",
  1478 => x"58a6f0c0",
  1479 => x"81c4496e",
  1480 => x"66dc4d69",
  1481 => x"a866d848",
  1482 => x"87c8c002",
  1483 => x"c048a6d8",
  1484 => x"87c5c078",
  1485 => x"c148a6d8",
  1486 => x"1e66d878",
  1487 => x"751ee0c0",
  1488 => x"d6deff49",
  1489 => x"7086c887",
  1490 => x"acb7c04c",
  1491 => x"87d4c106",
  1492 => x"e0c08574",
  1493 => x"75897449",
  1494 => x"dee1c14b",
  1495 => x"e5fe714a",
  1496 => x"85c287c6",
  1497 => x"4866e8c0",
  1498 => x"ecc080c1",
  1499 => x"ecc058a6",
  1500 => x"81c14966",
  1501 => x"c002a970",
  1502 => x"a6d887c8",
  1503 => x"c078c048",
  1504 => x"a6d887c5",
  1505 => x"d878c148",
  1506 => x"a4c21e66",
  1507 => x"48e0c049",
  1508 => x"49708871",
  1509 => x"ff49751e",
  1510 => x"c887c0dd",
  1511 => x"a8b7c086",
  1512 => x"87c0ff01",
  1513 => x"0266e8c0",
  1514 => x"6e87d1c0",
  1515 => x"c081c949",
  1516 => x"6e5166e8",
  1517 => x"efccc148",
  1518 => x"87ccc078",
  1519 => x"81c9496e",
  1520 => x"486e51c2",
  1521 => x"78e3cdc1",
  1522 => x"c6c07ec1",
  1523 => x"f6dbff87",
  1524 => x"6e4c7087",
  1525 => x"87f5c002",
  1526 => x"c84866c4",
  1527 => x"c004a866",
  1528 => x"66c487cb",
  1529 => x"c880c148",
  1530 => x"e0c058a6",
  1531 => x"4866c887",
  1532 => x"a6cc88c1",
  1533 => x"87d5c058",
  1534 => x"05acc6c1",
  1535 => x"cc87c8c0",
  1536 => x"80c14866",
  1537 => x"ff58a6d0",
  1538 => x"7087fcda",
  1539 => x"4866d04c",
  1540 => x"a6d480c1",
  1541 => x"029c7458",
  1542 => x"c487cbc0",
  1543 => x"c8c14866",
  1544 => x"f204a866",
  1545 => x"daff87ff",
  1546 => x"66c487d4",
  1547 => x"03a8c748",
  1548 => x"c387e5c0",
  1549 => x"c048d4c5",
  1550 => x"4966c478",
  1551 => x"c0c191cb",
  1552 => x"a1c48166",
  1553 => x"c04a6a4a",
  1554 => x"66c47952",
  1555 => x"c880c148",
  1556 => x"a8c758a6",
  1557 => x"87dbff04",
  1558 => x"e08ed0ff",
  1559 => x"203a87fb",
  1560 => x"1e731e00",
  1561 => x"029b4b71",
  1562 => x"c5c387c6",
  1563 => x"78c048d0",
  1564 => x"c5c31ec7",
  1565 => x"1e49bfd0",
  1566 => x"1ef7e4c1",
  1567 => x"bfccc5c3",
  1568 => x"87f4ee49",
  1569 => x"c5c386cc",
  1570 => x"e949bfcc",
  1571 => x"9b7387f9",
  1572 => x"c187c802",
  1573 => x"c049f7e4",
  1574 => x"ff87fce4",
  1575 => x"1e87fedf",
  1576 => x"c187d6c7",
  1577 => x"87f9fe49",
  1578 => x"87f4e9fe",
  1579 => x"cd029870",
  1580 => x"f1f2fe87",
  1581 => x"02987087",
  1582 => x"4ac187c4",
  1583 => x"4ac087c2",
  1584 => x"ce059a72",
  1585 => x"c11ec087",
  1586 => x"c049f0e3",
  1587 => x"c487fff2",
  1588 => x"c087fe86",
  1589 => x"fbe3c11e",
  1590 => x"f1f2c049",
  1591 => x"c11ec087",
  1592 => x"7087c8cf",
  1593 => x"e5f2c049",
  1594 => x"87ccc387",
  1595 => x"4f268ef8",
  1596 => x"66204453",
  1597 => x"656c6961",
  1598 => x"42002e64",
  1599 => x"69746f6f",
  1600 => x"2e2e676e",
  1601 => x"c01e002e",
  1602 => x"c087f0e7",
  1603 => x"f687caf6",
  1604 => x"1e4f2687",
  1605 => x"48d0c5c3",
  1606 => x"c5c378c0",
  1607 => x"78c048cc",
  1608 => x"e187fcfd",
  1609 => x"2648c087",
  1610 => x"4520804f",
  1611 => x"00746978",
  1612 => x"61422080",
  1613 => x"df006b63",
  1614 => x"65000012",
  1615 => x"00000031",
  1616 => x"12df0000",
  1617 => x"31830000",
  1618 => x"00000000",
  1619 => x"0012df00",
  1620 => x"0031a100",
  1621 => x"00000000",
  1622 => x"000012df",
  1623 => x"000031bf",
  1624 => x"df000000",
  1625 => x"dd000012",
  1626 => x"00000031",
  1627 => x"12df0000",
  1628 => x"31fb0000",
  1629 => x"00000000",
  1630 => x"0012df00",
  1631 => x"00321900",
  1632 => x"00000000",
  1633 => x"000012df",
  1634 => x"00000000",
  1635 => x"74000000",
  1636 => x"00000013",
  1637 => x"00000000",
  1638 => x"6f4c0000",
  1639 => x"2a206461",
  1640 => x"fe1e002e",
  1641 => x"78c048f0",
  1642 => x"097909cd",
  1643 => x"1e1e4f26",
  1644 => x"7ebff0fe",
  1645 => x"4f262648",
  1646 => x"48f0fe1e",
  1647 => x"4f2678c1",
  1648 => x"48f0fe1e",
  1649 => x"4f2678c0",
  1650 => x"c04a711e",
  1651 => x"4f265252",
  1652 => x"5c5b5e0e",
  1653 => x"86f40e5d",
  1654 => x"6d974d71",
  1655 => x"4ca5c17e",
  1656 => x"c8486c97",
  1657 => x"486e58a6",
  1658 => x"05a866c4",
  1659 => x"48ff87c5",
  1660 => x"ff87e6c0",
  1661 => x"a5c287ca",
  1662 => x"4b6c9749",
  1663 => x"974ba371",
  1664 => x"6c974b6b",
  1665 => x"c1486e7e",
  1666 => x"58a6c880",
  1667 => x"a6cc98c7",
  1668 => x"7c977058",
  1669 => x"7387e1fe",
  1670 => x"268ef448",
  1671 => x"264c264d",
  1672 => x"0e4f264b",
  1673 => x"0e5c5b5e",
  1674 => x"4c7186f4",
  1675 => x"c34a66d8",
  1676 => x"a4c29aff",
  1677 => x"496c974b",
  1678 => x"7249a173",
  1679 => x"7e6c9751",
  1680 => x"80c1486e",
  1681 => x"c758a6c8",
  1682 => x"58a6cc98",
  1683 => x"8ef45470",
  1684 => x"1e87caff",
  1685 => x"87e8fd1e",
  1686 => x"494abfe0",
  1687 => x"99c0e0c0",
  1688 => x"7287cb02",
  1689 => x"f7c8c31e",
  1690 => x"87f7fe49",
  1691 => x"fdfc86c4",
  1692 => x"fd7e7087",
  1693 => x"262687c2",
  1694 => x"c8c31e4f",
  1695 => x"c7fd49f7",
  1696 => x"d3e9c187",
  1697 => x"87dafc49",
  1698 => x"2687d0c5",
  1699 => x"5b5e0e4f",
  1700 => x"c30e5d5c",
  1701 => x"4abfd6c9",
  1702 => x"bfe1ebc1",
  1703 => x"bc724c49",
  1704 => x"dbfc4d71",
  1705 => x"744bc087",
  1706 => x"0299d049",
  1707 => x"497587d5",
  1708 => x"1e7199d0",
  1709 => x"f1c11ec0",
  1710 => x"82734aea",
  1711 => x"e4c04912",
  1712 => x"c186c887",
  1713 => x"c8832d2c",
  1714 => x"daff04ab",
  1715 => x"87e8fb87",
  1716 => x"48e1ebc1",
  1717 => x"bfd6c9c3",
  1718 => x"264d2678",
  1719 => x"264b264c",
  1720 => x"0000004f",
  1721 => x"d0ff1e00",
  1722 => x"78e1c848",
  1723 => x"c548d4ff",
  1724 => x"0266c478",
  1725 => x"e0c387c3",
  1726 => x"0266c878",
  1727 => x"d4ff87c6",
  1728 => x"78f0c348",
  1729 => x"7148d4ff",
  1730 => x"48d0ff78",
  1731 => x"c078e1c8",
  1732 => x"4f2678e0",
  1733 => x"5c5b5e0e",
  1734 => x"c34c710e",
  1735 => x"fa49f7c8",
  1736 => x"4a7087ee",
  1737 => x"04aab7c0",
  1738 => x"c387e3c2",
  1739 => x"c905aae0",
  1740 => x"d7efc187",
  1741 => x"c278c148",
  1742 => x"f0c387d4",
  1743 => x"87c905aa",
  1744 => x"48d3efc1",
  1745 => x"f5c178c1",
  1746 => x"d7efc187",
  1747 => x"87c702bf",
  1748 => x"c0c24b72",
  1749 => x"7287c2b3",
  1750 => x"059c744b",
  1751 => x"efc187d1",
  1752 => x"c11ebfd3",
  1753 => x"1ebfd7ef",
  1754 => x"f8fd4972",
  1755 => x"c186c887",
  1756 => x"02bfd3ef",
  1757 => x"7387e0c0",
  1758 => x"29b7c449",
  1759 => x"eaf0c191",
  1760 => x"cf4a7381",
  1761 => x"c192c29a",
  1762 => x"70307248",
  1763 => x"72baff4a",
  1764 => x"70986948",
  1765 => x"7387db79",
  1766 => x"29b7c449",
  1767 => x"eaf0c191",
  1768 => x"cf4a7381",
  1769 => x"c392c29a",
  1770 => x"70307248",
  1771 => x"b069484a",
  1772 => x"efc17970",
  1773 => x"78c048d7",
  1774 => x"48d3efc1",
  1775 => x"c8c378c0",
  1776 => x"cbf849f7",
  1777 => x"c04a7087",
  1778 => x"fd03aab7",
  1779 => x"48c087dd",
  1780 => x"0087c8fc",
  1781 => x"00000000",
  1782 => x"1e000000",
  1783 => x"49724ac0",
  1784 => x"f0c191c4",
  1785 => x"79c081ea",
  1786 => x"b7d082c1",
  1787 => x"87ee04aa",
  1788 => x"5e0e4f26",
  1789 => x"0e5d5c5b",
  1790 => x"c3f74d71",
  1791 => x"c44a7587",
  1792 => x"c1922ab7",
  1793 => x"7582eaf0",
  1794 => x"c29ccf4c",
  1795 => x"4b496a94",
  1796 => x"9bc32b74",
  1797 => x"307448c2",
  1798 => x"bcff4c70",
  1799 => x"98714874",
  1800 => x"d3f67a70",
  1801 => x"fa487387",
  1802 => x"000087ef",
  1803 => x"00000000",
  1804 => x"00000000",
  1805 => x"00000000",
  1806 => x"00000000",
  1807 => x"00000000",
  1808 => x"00000000",
  1809 => x"00000000",
  1810 => x"00000000",
  1811 => x"00000000",
  1812 => x"00000000",
  1813 => x"00000000",
  1814 => x"00000000",
  1815 => x"00000000",
  1816 => x"00000000",
  1817 => x"00000000",
  1818 => x"1e160000",
  1819 => x"362e2526",
  1820 => x"ff1e3e3d",
  1821 => x"e1c848d0",
  1822 => x"ff487178",
  1823 => x"267808d4",
  1824 => x"d0ff1e4f",
  1825 => x"78e1c848",
  1826 => x"d4ff4871",
  1827 => x"66c47808",
  1828 => x"08d4ff48",
  1829 => x"1e4f2678",
  1830 => x"66c44a71",
  1831 => x"49721e49",
  1832 => x"ff87deff",
  1833 => x"e0c048d0",
  1834 => x"4f262678",
  1835 => x"c24a711e",
  1836 => x"c303aab7",
  1837 => x"87c28287",
  1838 => x"66c482ce",
  1839 => x"ff49721e",
  1840 => x"262687d5",
  1841 => x"d4ff1e4f",
  1842 => x"7affc34a",
  1843 => x"c848d0ff",
  1844 => x"7ade78e1",
  1845 => x"bfc1c9c3",
  1846 => x"c848497a",
  1847 => x"717a7028",
  1848 => x"7028d048",
  1849 => x"d848717a",
  1850 => x"ff7a7028",
  1851 => x"e0c048d0",
  1852 => x"0e4f2678",
  1853 => x"5d5c5b5e",
  1854 => x"c34c710e",
  1855 => x"4dbfc1c9",
  1856 => x"d02b744b",
  1857 => x"83c19b66",
  1858 => x"04ab66d4",
  1859 => x"4bc087c2",
  1860 => x"66d04a74",
  1861 => x"ff317249",
  1862 => x"739975b9",
  1863 => x"70307248",
  1864 => x"b071484a",
  1865 => x"58c5c9c3",
  1866 => x"2687dafe",
  1867 => x"264c264d",
  1868 => x"1e4f264b",
  1869 => x"c848d0ff",
  1870 => x"487178c9",
  1871 => x"7808d4ff",
  1872 => x"711e4f26",
  1873 => x"87eb494a",
  1874 => x"c848d0ff",
  1875 => x"1e4f2678",
  1876 => x"4b711e73",
  1877 => x"bfd1c9c3",
  1878 => x"c287c302",
  1879 => x"d0ff87eb",
  1880 => x"78c9c848",
  1881 => x"e0c04973",
  1882 => x"48d4ffb1",
  1883 => x"c9c37871",
  1884 => x"78c048c5",
  1885 => x"c50266c8",
  1886 => x"49ffc387",
  1887 => x"49c087c2",
  1888 => x"59cdc9c3",
  1889 => x"c60266cc",
  1890 => x"d5d5c587",
  1891 => x"cf87c44a",
  1892 => x"c34affff",
  1893 => x"c35ad1c9",
  1894 => x"c148d1c9",
  1895 => x"2687c478",
  1896 => x"264c264d",
  1897 => x"0e4f264b",
  1898 => x"5d5c5b5e",
  1899 => x"c34a710e",
  1900 => x"4cbfcdc9",
  1901 => x"cb029a72",
  1902 => x"91c84987",
  1903 => x"4bc5f5c1",
  1904 => x"87c48371",
  1905 => x"4bc5f9c1",
  1906 => x"49134dc0",
  1907 => x"c9c39974",
  1908 => x"ffb9bfc9",
  1909 => x"787148d4",
  1910 => x"852cb7c1",
  1911 => x"04adb7c8",
  1912 => x"c9c387e8",
  1913 => x"c848bfc5",
  1914 => x"c9c9c380",
  1915 => x"87effe58",
  1916 => x"711e731e",
  1917 => x"9a4a134b",
  1918 => x"7287cb02",
  1919 => x"87e7fe49",
  1920 => x"059a4a13",
  1921 => x"dafe87f5",
  1922 => x"c9c31e87",
  1923 => x"c349bfc5",
  1924 => x"c148c5c9",
  1925 => x"c0c478a1",
  1926 => x"db03a9b7",
  1927 => x"48d4ff87",
  1928 => x"bfc9c9c3",
  1929 => x"c5c9c378",
  1930 => x"c9c349bf",
  1931 => x"a1c148c5",
  1932 => x"b7c0c478",
  1933 => x"87e504a9",
  1934 => x"c848d0ff",
  1935 => x"d1c9c378",
  1936 => x"2678c048",
  1937 => x"0000004f",
  1938 => x"00000000",
  1939 => x"00000000",
  1940 => x"00005f5f",
  1941 => x"03030000",
  1942 => x"00030300",
  1943 => x"7f7f1400",
  1944 => x"147f7f14",
  1945 => x"2e240000",
  1946 => x"123a6b6b",
  1947 => x"366a4c00",
  1948 => x"32566c18",
  1949 => x"4f7e3000",
  1950 => x"683a7759",
  1951 => x"04000040",
  1952 => x"00000307",
  1953 => x"1c000000",
  1954 => x"0041633e",
  1955 => x"41000000",
  1956 => x"001c3e63",
  1957 => x"3e2a0800",
  1958 => x"2a3e1c1c",
  1959 => x"08080008",
  1960 => x"08083e3e",
  1961 => x"80000000",
  1962 => x"000060e0",
  1963 => x"08080000",
  1964 => x"08080808",
  1965 => x"00000000",
  1966 => x"00006060",
  1967 => x"30604000",
  1968 => x"03060c18",
  1969 => x"7f3e0001",
  1970 => x"3e7f4d59",
  1971 => x"06040000",
  1972 => x"00007f7f",
  1973 => x"63420000",
  1974 => x"464f5971",
  1975 => x"63220000",
  1976 => x"367f4949",
  1977 => x"161c1800",
  1978 => x"107f7f13",
  1979 => x"67270000",
  1980 => x"397d4545",
  1981 => x"7e3c0000",
  1982 => x"3079494b",
  1983 => x"01010000",
  1984 => x"070f7971",
  1985 => x"7f360000",
  1986 => x"367f4949",
  1987 => x"4f060000",
  1988 => x"1e3f6949",
  1989 => x"00000000",
  1990 => x"00006666",
  1991 => x"80000000",
  1992 => x"000066e6",
  1993 => x"08080000",
  1994 => x"22221414",
  1995 => x"14140000",
  1996 => x"14141414",
  1997 => x"22220000",
  1998 => x"08081414",
  1999 => x"03020000",
  2000 => x"060f5951",
  2001 => x"417f3e00",
  2002 => x"1e1f555d",
  2003 => x"7f7e0000",
  2004 => x"7e7f0909",
  2005 => x"7f7f0000",
  2006 => x"367f4949",
  2007 => x"3e1c0000",
  2008 => x"41414163",
  2009 => x"7f7f0000",
  2010 => x"1c3e6341",
  2011 => x"7f7f0000",
  2012 => x"41414949",
  2013 => x"7f7f0000",
  2014 => x"01010909",
  2015 => x"7f3e0000",
  2016 => x"7a7b4941",
  2017 => x"7f7f0000",
  2018 => x"7f7f0808",
  2019 => x"41000000",
  2020 => x"00417f7f",
  2021 => x"60200000",
  2022 => x"3f7f4040",
  2023 => x"087f7f00",
  2024 => x"4163361c",
  2025 => x"7f7f0000",
  2026 => x"40404040",
  2027 => x"067f7f00",
  2028 => x"7f7f060c",
  2029 => x"067f7f00",
  2030 => x"7f7f180c",
  2031 => x"7f3e0000",
  2032 => x"3e7f4141",
  2033 => x"7f7f0000",
  2034 => x"060f0909",
  2035 => x"417f3e00",
  2036 => x"407e7f61",
  2037 => x"7f7f0000",
  2038 => x"667f1909",
  2039 => x"6f260000",
  2040 => x"327b594d",
  2041 => x"01010000",
  2042 => x"01017f7f",
  2043 => x"7f3f0000",
  2044 => x"3f7f4040",
  2045 => x"3f0f0000",
  2046 => x"0f3f7070",
  2047 => x"307f7f00",
  2048 => x"7f7f3018",
  2049 => x"36634100",
  2050 => x"63361c1c",
  2051 => x"06030141",
  2052 => x"03067c7c",
  2053 => x"59716101",
  2054 => x"4143474d",
  2055 => x"7f000000",
  2056 => x"0041417f",
  2057 => x"06030100",
  2058 => x"6030180c",
  2059 => x"41000040",
  2060 => x"007f7f41",
  2061 => x"060c0800",
  2062 => x"080c0603",
  2063 => x"80808000",
  2064 => x"80808080",
  2065 => x"00000000",
  2066 => x"00040703",
  2067 => x"74200000",
  2068 => x"787c5454",
  2069 => x"7f7f0000",
  2070 => x"387c4444",
  2071 => x"7c380000",
  2072 => x"00444444",
  2073 => x"7c380000",
  2074 => x"7f7f4444",
  2075 => x"7c380000",
  2076 => x"185c5454",
  2077 => x"7e040000",
  2078 => x"0005057f",
  2079 => x"bc180000",
  2080 => x"7cfca4a4",
  2081 => x"7f7f0000",
  2082 => x"787c0404",
  2083 => x"00000000",
  2084 => x"00407d3d",
  2085 => x"80800000",
  2086 => x"007dfd80",
  2087 => x"7f7f0000",
  2088 => x"446c3810",
  2089 => x"00000000",
  2090 => x"00407f3f",
  2091 => x"0c7c7c00",
  2092 => x"787c0c18",
  2093 => x"7c7c0000",
  2094 => x"787c0404",
  2095 => x"7c380000",
  2096 => x"387c4444",
  2097 => x"fcfc0000",
  2098 => x"183c2424",
  2099 => x"3c180000",
  2100 => x"fcfc2424",
  2101 => x"7c7c0000",
  2102 => x"080c0404",
  2103 => x"5c480000",
  2104 => x"20745454",
  2105 => x"3f040000",
  2106 => x"0044447f",
  2107 => x"7c3c0000",
  2108 => x"7c7c4040",
  2109 => x"3c1c0000",
  2110 => x"1c3c6060",
  2111 => x"607c3c00",
  2112 => x"3c7c6030",
  2113 => x"386c4400",
  2114 => x"446c3810",
  2115 => x"bc1c0000",
  2116 => x"1c3c60e0",
  2117 => x"64440000",
  2118 => x"444c5c74",
  2119 => x"08080000",
  2120 => x"4141773e",
  2121 => x"00000000",
  2122 => x"00007f7f",
  2123 => x"41410000",
  2124 => x"08083e77",
  2125 => x"01010200",
  2126 => x"01020203",
  2127 => x"7f7f7f00",
  2128 => x"7f7f7f7f",
  2129 => x"1c080800",
  2130 => x"7f3e3e1c",
  2131 => x"3e7f7f7f",
  2132 => x"081c1c3e",
  2133 => x"18100008",
  2134 => x"10187c7c",
  2135 => x"30100000",
  2136 => x"10307c7c",
  2137 => x"60301000",
  2138 => x"061e7860",
  2139 => x"3c664200",
  2140 => x"42663c18",
  2141 => x"6a387800",
  2142 => x"386cc6c2",
  2143 => x"00006000",
  2144 => x"60000060",
  2145 => x"5b5e0e00",
  2146 => x"1e0e5d5c",
  2147 => x"c9c34c71",
  2148 => x"c04dbfe2",
  2149 => x"741ec04b",
  2150 => x"87c702ab",
  2151 => x"c048a6c4",
  2152 => x"c487c578",
  2153 => x"78c148a6",
  2154 => x"731e66c4",
  2155 => x"87dfee49",
  2156 => x"e0c086c8",
  2157 => x"87efef49",
  2158 => x"6a4aa5c4",
  2159 => x"87f0f049",
  2160 => x"cb87c6f1",
  2161 => x"c883c185",
  2162 => x"ff04abb7",
  2163 => x"262687c7",
  2164 => x"264c264d",
  2165 => x"1e4f264b",
  2166 => x"c9c34a71",
  2167 => x"c9c35ae6",
  2168 => x"78c748e6",
  2169 => x"87ddfe49",
  2170 => x"731e4f26",
  2171 => x"c04a711e",
  2172 => x"d303aab7",
  2173 => x"f8d7c287",
  2174 => x"87c405bf",
  2175 => x"87c24bc1",
  2176 => x"d7c24bc0",
  2177 => x"87c45bfc",
  2178 => x"5afcd7c2",
  2179 => x"bff8d7c2",
  2180 => x"c19ac14a",
  2181 => x"ec49a2c0",
  2182 => x"d7c287e8",
  2183 => x"c249bfe0",
  2184 => x"b1bff8d7",
  2185 => x"787148fc",
  2186 => x"1e87e8fe",
  2187 => x"66c44a71",
  2188 => x"e949721e",
  2189 => x"262687f6",
  2190 => x"d7c21e4f",
  2191 => x"c049bff8",
  2192 => x"c387d7e9",
  2193 => x"e848dac9",
  2194 => x"c9c378bf",
  2195 => x"bfec48d6",
  2196 => x"dac9c378",
  2197 => x"c3494abf",
  2198 => x"b7c899ff",
  2199 => x"7148722a",
  2200 => x"e2c9c3b0",
  2201 => x"0e4f2658",
  2202 => x"5d5c5b5e",
  2203 => x"ff4b710e",
  2204 => x"c9c387c7",
  2205 => x"50c048d5",
  2206 => x"f5e54973",
  2207 => x"4c497087",
  2208 => x"eecb9cc2",
  2209 => x"87f8cd49",
  2210 => x"c34d4970",
  2211 => x"bf97d5c9",
  2212 => x"87e2c105",
  2213 => x"c34966d0",
  2214 => x"99bfdec9",
  2215 => x"d487d605",
  2216 => x"c9c34966",
  2217 => x"0599bfd6",
  2218 => x"497387cb",
  2219 => x"7087c3e5",
  2220 => x"c1c10298",
  2221 => x"fd4cc187",
  2222 => x"497587ff",
  2223 => x"7087cdcd",
  2224 => x"87c60298",
  2225 => x"48d5c9c3",
  2226 => x"c9c350c1",
  2227 => x"05bf97d5",
  2228 => x"c387e3c0",
  2229 => x"49bfdec9",
  2230 => x"059966d0",
  2231 => x"c387d6ff",
  2232 => x"49bfd6c9",
  2233 => x"059966d4",
  2234 => x"7387caff",
  2235 => x"87c2e449",
  2236 => x"fe059870",
  2237 => x"487487ff",
  2238 => x"0e87d4fb",
  2239 => x"5d5c5b5e",
  2240 => x"c086f80e",
  2241 => x"bfec4c4d",
  2242 => x"48a6c47e",
  2243 => x"bfe2c9c3",
  2244 => x"1e1ec078",
  2245 => x"fd49f7c1",
  2246 => x"86c887cd",
  2247 => x"c0029870",
  2248 => x"d7c287f3",
  2249 => x"c405bfe0",
  2250 => x"c27ec187",
  2251 => x"c27ec087",
  2252 => x"6e48e0d7",
  2253 => x"1efcca78",
  2254 => x"c90266c4",
  2255 => x"48a6c487",
  2256 => x"78f7d5c2",
  2257 => x"a6c487c7",
  2258 => x"c2d6c248",
  2259 => x"4966c478",
  2260 => x"c487fbc8",
  2261 => x"c01ec186",
  2262 => x"fc49c71e",
  2263 => x"86c887c9",
  2264 => x"cd029870",
  2265 => x"fa49ff87",
  2266 => x"dac187c0",
  2267 => x"87c2e249",
  2268 => x"c9c34dc1",
  2269 => x"02bf97d5",
  2270 => x"f4d687c3",
  2271 => x"dac9c387",
  2272 => x"d7c24bbf",
  2273 => x"c105bff8",
  2274 => x"d7c287e1",
  2275 => x"c002bfe0",
  2276 => x"a6c487f0",
  2277 => x"c0c0c848",
  2278 => x"e4d7c278",
  2279 => x"bf976e7e",
  2280 => x"c1486e49",
  2281 => x"717e7080",
  2282 => x"7087c7e1",
  2283 => x"87c30298",
  2284 => x"c4b366c4",
  2285 => x"b7c14866",
  2286 => x"58a6c828",
  2287 => x"ff059870",
  2288 => x"fdc387db",
  2289 => x"87eae049",
  2290 => x"e049fac3",
  2291 => x"497387e4",
  2292 => x"7199ffc3",
  2293 => x"f949c01e",
  2294 => x"497387d1",
  2295 => x"7129b7c8",
  2296 => x"f949c11e",
  2297 => x"86c887c5",
  2298 => x"c387c7c6",
  2299 => x"4bbfdec9",
  2300 => x"87df029b",
  2301 => x"bff4d7c2",
  2302 => x"87d0c849",
  2303 => x"c0059870",
  2304 => x"4bc087c4",
  2305 => x"e0c287d3",
  2306 => x"87f4c749",
  2307 => x"58f8d7c2",
  2308 => x"c287c6c0",
  2309 => x"c048f4d7",
  2310 => x"c2497378",
  2311 => x"cfc00599",
  2312 => x"49ebc387",
  2313 => x"87cadfff",
  2314 => x"99c24970",
  2315 => x"87c2c002",
  2316 => x"49734cfb",
  2317 => x"c00599c1",
  2318 => x"f4c387cf",
  2319 => x"f1deff49",
  2320 => x"c2497087",
  2321 => x"c2c00299",
  2322 => x"734cfa87",
  2323 => x"0599c849",
  2324 => x"c387cfc0",
  2325 => x"deff49f5",
  2326 => x"497087d8",
  2327 => x"c00299c2",
  2328 => x"c9c387d6",
  2329 => x"c002bfe6",
  2330 => x"c14887ca",
  2331 => x"eac9c388",
  2332 => x"87c2c058",
  2333 => x"4dc14cff",
  2334 => x"99c44973",
  2335 => x"87cfc005",
  2336 => x"ff49f2c3",
  2337 => x"7087ebdd",
  2338 => x"0299c249",
  2339 => x"c387dcc0",
  2340 => x"7ebfe6c9",
  2341 => x"a8b7c748",
  2342 => x"87cbc003",
  2343 => x"80c1486e",
  2344 => x"58eac9c3",
  2345 => x"fe87c2c0",
  2346 => x"c34dc14c",
  2347 => x"ddff49fd",
  2348 => x"497087c0",
  2349 => x"c00299c2",
  2350 => x"c9c387d5",
  2351 => x"c002bfe6",
  2352 => x"c9c387c9",
  2353 => x"78c048e6",
  2354 => x"fd87c2c0",
  2355 => x"c34dc14c",
  2356 => x"dcff49fa",
  2357 => x"497087dc",
  2358 => x"c00299c2",
  2359 => x"c9c387d9",
  2360 => x"c748bfe6",
  2361 => x"c003a8b7",
  2362 => x"c9c387c9",
  2363 => x"78c748e6",
  2364 => x"fc87c2c0",
  2365 => x"c04dc14c",
  2366 => x"c003acb7",
  2367 => x"66c487d5",
  2368 => x"80d8c148",
  2369 => x"bf6e7e70",
  2370 => x"87c7c002",
  2371 => x"744bbf6e",
  2372 => x"c00f7349",
  2373 => x"1ef0c31e",
  2374 => x"f549dac1",
  2375 => x"86c887c9",
  2376 => x"c0029870",
  2377 => x"c9c387d9",
  2378 => x"6e7ebfe6",
  2379 => x"c491cb49",
  2380 => x"82714a66",
  2381 => x"c6c0026a",
  2382 => x"6e4b6a87",
  2383 => x"750f7349",
  2384 => x"c8c0029d",
  2385 => x"e6c9c387",
  2386 => x"f8f049bf",
  2387 => x"fcd7c287",
  2388 => x"ddc002bf",
  2389 => x"f3c24987",
  2390 => x"02987087",
  2391 => x"c387d3c0",
  2392 => x"49bfe6c9",
  2393 => x"c087def0",
  2394 => x"87fef149",
  2395 => x"48fcd7c2",
  2396 => x"8ef878c0",
  2397 => x"4a87d8f1",
  2398 => x"656b796f",
  2399 => x"6f207379",
  2400 => x"6f4a006e",
  2401 => x"79656b79",
  2402 => x"666f2073",
  2403 => x"5e0e0066",
  2404 => x"0e5d5c5b",
  2405 => x"c34c711e",
  2406 => x"49bfe2c9",
  2407 => x"4da1cdc1",
  2408 => x"6981d1c1",
  2409 => x"029c747e",
  2410 => x"a5c487cf",
  2411 => x"c37b744b",
  2412 => x"49bfe2c9",
  2413 => x"6e87e0f0",
  2414 => x"059c747b",
  2415 => x"4bc087c4",
  2416 => x"4bc187c2",
  2417 => x"e1f04973",
  2418 => x"0266d487",
  2419 => x"c04987c8",
  2420 => x"4a7087ee",
  2421 => x"4ac087c2",
  2422 => x"5ac0d8c2",
  2423 => x"87efef26",
  2424 => x"00000000",
  2425 => x"14111258",
  2426 => x"231c1b1d",
  2427 => x"9491595a",
  2428 => x"f4ebf2f5",
  2429 => x"00000000",
  2430 => x"00000000",
  2431 => x"00000000",
  2432 => x"ff4a711e",
  2433 => x"7249bfc8",
  2434 => x"4f2648a1",
  2435 => x"bfc8ff1e",
  2436 => x"c0c0fe89",
  2437 => x"a9c0c0c0",
  2438 => x"c087c401",
  2439 => x"c187c24a",
  2440 => x"2648724a",
  2441 => x"5b5e0e4f",
  2442 => x"710e5d5c",
  2443 => x"4cd4ff4b",
  2444 => x"c04866d0",
  2445 => x"ff49d678",
  2446 => x"c387f7d8",
  2447 => x"496c7cff",
  2448 => x"7199ffc3",
  2449 => x"f0c3494d",
  2450 => x"a9e0c199",
  2451 => x"c387cb05",
  2452 => x"486c7cff",
  2453 => x"66d098c3",
  2454 => x"ffc37808",
  2455 => x"494a6c7c",
  2456 => x"ffc331c8",
  2457 => x"714a6c7c",
  2458 => x"c84972b2",
  2459 => x"7cffc331",
  2460 => x"b2714a6c",
  2461 => x"31c84972",
  2462 => x"6c7cffc3",
  2463 => x"ffb2714a",
  2464 => x"e0c048d0",
  2465 => x"029b7378",
  2466 => x"7b7287c2",
  2467 => x"4d264875",
  2468 => x"4b264c26",
  2469 => x"261e4f26",
  2470 => x"5b5e0e4f",
  2471 => x"86f80e5c",
  2472 => x"a6c81e76",
  2473 => x"87fdfd49",
  2474 => x"4b7086c4",
  2475 => x"a8c2486e",
  2476 => x"87cac303",
  2477 => x"f0c34a73",
  2478 => x"aad0c19a",
  2479 => x"c187c702",
  2480 => x"c205aae0",
  2481 => x"497387f8",
  2482 => x"c30299c8",
  2483 => x"87c6ff87",
  2484 => x"9cc34c73",
  2485 => x"c105acc2",
  2486 => x"66c487cf",
  2487 => x"7131c949",
  2488 => x"4a66c41e",
  2489 => x"c392c8c1",
  2490 => x"7249eac9",
  2491 => x"ded0fe81",
  2492 => x"4966c487",
  2493 => x"49e3c01e",
  2494 => x"87dbd6ff",
  2495 => x"d5ff49d8",
  2496 => x"c0c887f0",
  2497 => x"daf8c21e",
  2498 => x"f3e8fd49",
  2499 => x"48d0ff87",
  2500 => x"c278e0c0",
  2501 => x"d01edaf8",
  2502 => x"c8c14a66",
  2503 => x"eac9c392",
  2504 => x"fe817249",
  2505 => x"d087e6cb",
  2506 => x"05acc186",
  2507 => x"c487cfc1",
  2508 => x"31c94966",
  2509 => x"66c41e71",
  2510 => x"92c8c14a",
  2511 => x"49eac9c3",
  2512 => x"cffe8172",
  2513 => x"f8c287c9",
  2514 => x"66c81eda",
  2515 => x"92c8c14a",
  2516 => x"49eac9c3",
  2517 => x"c9fe8172",
  2518 => x"66c887f0",
  2519 => x"e3c01e49",
  2520 => x"f2d4ff49",
  2521 => x"ff49d787",
  2522 => x"c887c7d4",
  2523 => x"f8c21ec0",
  2524 => x"e6fd49da",
  2525 => x"86d087f4",
  2526 => x"c048d0ff",
  2527 => x"8ef878e0",
  2528 => x"0e87cdfc",
  2529 => x"5d5c5b5e",
  2530 => x"4d711e0e",
  2531 => x"d44cd4ff",
  2532 => x"c3487e66",
  2533 => x"c506a8b7",
  2534 => x"c148c087",
  2535 => x"497587e3",
  2536 => x"87d2dffe",
  2537 => x"66c41e75",
  2538 => x"93c8c14b",
  2539 => x"83eac9c3",
  2540 => x"c3fe4973",
  2541 => x"83c887fe",
  2542 => x"d0ff4b6b",
  2543 => x"78e1c848",
  2544 => x"49737cdd",
  2545 => x"7199ffc3",
  2546 => x"c849737c",
  2547 => x"ffc329b7",
  2548 => x"737c7199",
  2549 => x"29b7d049",
  2550 => x"7199ffc3",
  2551 => x"d849737c",
  2552 => x"7c7129b7",
  2553 => x"7c7c7cc0",
  2554 => x"7c7c7c7c",
  2555 => x"7c7c7c7c",
  2556 => x"78e0c07c",
  2557 => x"dc1e66c4",
  2558 => x"dad2ff49",
  2559 => x"7386c887",
  2560 => x"c9fa2648",
  2561 => x"5b5e0e87",
  2562 => x"1e0e5d5c",
  2563 => x"d4ff7e71",
  2564 => x"c31e6e4b",
  2565 => x"fe49facb",
  2566 => x"c487d9c2",
  2567 => x"9d4d7086",
  2568 => x"87c3c302",
  2569 => x"bfc2ccc3",
  2570 => x"fe496e4c",
  2571 => x"ff87c7dd",
  2572 => x"c5c848d0",
  2573 => x"7bd6c178",
  2574 => x"7b154ac0",
  2575 => x"e0c082c1",
  2576 => x"f504aab7",
  2577 => x"48d0ff87",
  2578 => x"c5c878c4",
  2579 => x"7bd3c178",
  2580 => x"78c47bc1",
  2581 => x"c1029c74",
  2582 => x"f8c287fc",
  2583 => x"c0c87eda",
  2584 => x"b7c08c4d",
  2585 => x"87c603ac",
  2586 => x"4da4c0c8",
  2587 => x"c5c34cc0",
  2588 => x"49bf97cb",
  2589 => x"d20299d0",
  2590 => x"c31ec087",
  2591 => x"fe49facb",
  2592 => x"c487c7c5",
  2593 => x"4a497086",
  2594 => x"c287efc0",
  2595 => x"c31edaf8",
  2596 => x"fe49facb",
  2597 => x"c487f3c4",
  2598 => x"4a497086",
  2599 => x"c848d0ff",
  2600 => x"d4c178c5",
  2601 => x"bf976e7b",
  2602 => x"c1486e7b",
  2603 => x"c17e7080",
  2604 => x"f0ff058d",
  2605 => x"48d0ff87",
  2606 => x"9a7278c4",
  2607 => x"c087c505",
  2608 => x"87e5c048",
  2609 => x"cbc31ec1",
  2610 => x"c2fe49fa",
  2611 => x"86c487db",
  2612 => x"fe059c74",
  2613 => x"d0ff87c4",
  2614 => x"78c5c848",
  2615 => x"c07bd3c1",
  2616 => x"c178c47b",
  2617 => x"c087c248",
  2618 => x"4d262648",
  2619 => x"4b264c26",
  2620 => x"5e0e4f26",
  2621 => x"710e5c5b",
  2622 => x"0266cc4b",
  2623 => x"c04c87d8",
  2624 => x"d8028cf0",
  2625 => x"c14a7487",
  2626 => x"87d1028a",
  2627 => x"87cd028a",
  2628 => x"87c9028a",
  2629 => x"497387d7",
  2630 => x"d087eafb",
  2631 => x"c01e7487",
  2632 => x"87dff949",
  2633 => x"49731e74",
  2634 => x"c887d8f9",
  2635 => x"87fcfe86",
  2636 => x"e5c21e00",
  2637 => x"c149bfda",
  2638 => x"dee5c2b9",
  2639 => x"48d4ff59",
  2640 => x"ff78ffc3",
  2641 => x"e1c848d0",
  2642 => x"48d4ff78",
  2643 => x"31c478c1",
  2644 => x"d0ff7871",
  2645 => x"78e0c048",
  2646 => x"00004f26",
  2647 => x"ff1e0000",
  2648 => x"c487ddc1",
  2649 => x"c0c24966",
  2650 => x"87cd0299",
  2651 => x"c31ee0c3",
  2652 => x"ff49f7c8",
  2653 => x"c487ecc2",
  2654 => x"4966c486",
  2655 => x"0299c0c4",
  2656 => x"f0c387cd",
  2657 => x"f7c8c31e",
  2658 => x"d6c2ff49",
  2659 => x"c486c487",
  2660 => x"ffc14966",
  2661 => x"c31e7199",
  2662 => x"ff49f7c8",
  2663 => x"ff87c4c2",
  2664 => x"2687d5c0",
  2665 => x"5e0e4f26",
  2666 => x"0e5d5c5b",
  2667 => x"c086d8ff",
  2668 => x"c6cdc37e",
  2669 => x"81c249bf",
  2670 => x"1e721e71",
  2671 => x"dcfd4ac6",
  2672 => x"487187f7",
  2673 => x"49264a26",
  2674 => x"c358a6c8",
  2675 => x"49bfc6cd",
  2676 => x"1e7181c4",
  2677 => x"4ac61e72",
  2678 => x"87dddcfd",
  2679 => x"4a264871",
  2680 => x"a6cc4926",
  2681 => x"f7f1c258",
  2682 => x"dff049bf",
  2683 => x"02987087",
  2684 => x"c087f9c9",
  2685 => x"c7f049e0",
  2686 => x"c2497087",
  2687 => x"c059fbf1",
  2688 => x"c449744c",
  2689 => x"81d0fe91",
  2690 => x"49744a69",
  2691 => x"bfc6cdc3",
  2692 => x"c391c481",
  2693 => x"7281d2cd",
  2694 => x"d2029a79",
  2695 => x"c1497287",
  2696 => x"6e9a7189",
  2697 => x"7080c148",
  2698 => x"059a727e",
  2699 => x"c187eeff",
  2700 => x"acb7c284",
  2701 => x"87c9ff04",
  2702 => x"fcc0486e",
  2703 => x"c804a8b7",
  2704 => x"4cc087ea",
  2705 => x"66c44a74",
  2706 => x"c392c482",
  2707 => x"7482d2cd",
  2708 => x"8166c849",
  2709 => x"cdc391c4",
  2710 => x"4a6a81d2",
  2711 => x"b9724969",
  2712 => x"cdc34b74",
  2713 => x"c483bfc6",
  2714 => x"d2cdc393",
  2715 => x"72ba6b83",
  2716 => x"d4987148",
  2717 => x"497458a6",
  2718 => x"bfc6cdc3",
  2719 => x"c391c481",
  2720 => x"6981d2cd",
  2721 => x"48a6d47e",
  2722 => x"a6d078c0",
  2723 => x"4cffc35c",
  2724 => x"df4966d0",
  2725 => x"e2c60229",
  2726 => x"4a66cc87",
  2727 => x"d492e0c0",
  2728 => x"ffc08266",
  2729 => x"70887248",
  2730 => x"48a6d84a",
  2731 => x"80c478c0",
  2732 => x"496e78c0",
  2733 => x"e4c029df",
  2734 => x"cdc359a6",
  2735 => x"78c148c2",
  2736 => x"31c34972",
  2737 => x"b1722ab7",
  2738 => x"c499ffc0",
  2739 => x"f3f3c291",
  2740 => x"6d85714d",
  2741 => x"c0c4494b",
  2742 => x"d70299c0",
  2743 => x"66e0c087",
  2744 => x"87c7c002",
  2745 => x"78c080c8",
  2746 => x"c387d0c5",
  2747 => x"c148cacd",
  2748 => x"87c7c578",
  2749 => x"0266e0c0",
  2750 => x"497387d8",
  2751 => x"99c0c0c2",
  2752 => x"87c3c002",
  2753 => x"6d2bb7d0",
  2754 => x"fffffd48",
  2755 => x"c07d7098",
  2756 => x"cdc387fa",
  2757 => x"c002bfca",
  2758 => x"487387f2",
  2759 => x"c028b7d0",
  2760 => x"7058a6e8",
  2761 => x"e3c00298",
  2762 => x"cecdc387",
  2763 => x"e0c049bf",
  2764 => x"c00299c0",
  2765 => x"497087ca",
  2766 => x"99c0e0c0",
  2767 => x"87ccc002",
  2768 => x"c0c2486d",
  2769 => x"7d70b0c0",
  2770 => x"4b66e4c0",
  2771 => x"c0c84973",
  2772 => x"c20299c0",
  2773 => x"cdc387c5",
  2774 => x"cc4abfce",
  2775 => x"c0029ac0",
  2776 => x"c0c487cf",
  2777 => x"d7c0028a",
  2778 => x"c0028a87",
  2779 => x"dcc187f8",
  2780 => x"74497387",
  2781 => x"c291c299",
  2782 => x"1181e7f3",
  2783 => x"87dbc14b",
  2784 => x"99744973",
  2785 => x"f3c291c2",
  2786 => x"81c181e7",
  2787 => x"e0c04b11",
  2788 => x"c8c00266",
  2789 => x"48a6dc87",
  2790 => x"fec078d2",
  2791 => x"48a6d887",
  2792 => x"c078d2c4",
  2793 => x"497387f5",
  2794 => x"91c29974",
  2795 => x"81e7f3c2",
  2796 => x"4b1181c1",
  2797 => x"0266e0c0",
  2798 => x"dc87c9c0",
  2799 => x"d9c148a6",
  2800 => x"87d7c078",
  2801 => x"c548a6d8",
  2802 => x"cec078d9",
  2803 => x"74497387",
  2804 => x"c291c299",
  2805 => x"c181e7f3",
  2806 => x"c04b1181",
  2807 => x"c00266e0",
  2808 => x"497387db",
  2809 => x"fcc7b9ff",
  2810 => x"487199c0",
  2811 => x"bfcecdc3",
  2812 => x"d2cdc398",
  2813 => x"c49b7458",
  2814 => x"d3c0b3c0",
  2815 => x"c7497387",
  2816 => x"7199c0fc",
  2817 => x"cecdc348",
  2818 => x"cdc3b0bf",
  2819 => x"9b7458d2",
  2820 => x"c00266d8",
  2821 => x"c31e87ca",
  2822 => x"f549c2cd",
  2823 => x"86c487c0",
  2824 => x"cdc31e73",
  2825 => x"f5f449c2",
  2826 => x"dc86c487",
  2827 => x"cac00266",
  2828 => x"cdc31e87",
  2829 => x"e5f449c2",
  2830 => x"d086c487",
  2831 => x"30c14866",
  2832 => x"6e58a6d4",
  2833 => x"7030c148",
  2834 => x"4866d47e",
  2835 => x"a6d880c1",
  2836 => x"b7e0c058",
  2837 => x"f7f804a8",
  2838 => x"4c66cc87",
  2839 => x"b7c284c1",
  2840 => x"dff704ac",
  2841 => x"c6cdc387",
  2842 => x"7866c448",
  2843 => x"268ed8ff",
  2844 => x"264c264d",
  2845 => x"004f264b",
  2846 => x"1e000000",
  2847 => x"49724ac0",
  2848 => x"cdc391c4",
  2849 => x"79ff81d2",
  2850 => x"b7c682c1",
  2851 => x"87ee04aa",
  2852 => x"48c6cdc3",
  2853 => x"784040c0",
  2854 => x"731e4f26",
  2855 => x"f44b711e",
  2856 => x"497387c4",
  2857 => x"87ecf9fe",
  2858 => x"1e87c8ff",
  2859 => x"4bc01e73",
  2860 => x"49c8f3c2",
  2861 => x"7087ceed",
  2862 => x"87c40598",
  2863 => x"4bd4f3c2",
  2864 => x"7387f8fe",
  2865 => x"87ebfe48",
  2866 => x"4349524f",
  2867 => x"20202020",
  2868 => x"004d4f52",
  2869 => x"204d4f52",
  2870 => x"64616f6c",
  2871 => x"20676e69",
  2872 => x"6c696166",
  2873 => x"f4006465",
  2874 => x"05f5f2eb",
  2875 => x"030c0406",
  2876 => x"660a830b",
  2877 => x"5a00fc00",
  2878 => x"0000da00",
  2879 => x"05089480",
  2880 => x"02007880",
  2881 => x"03000180",
  2882 => x"04000980",
  2883 => x"01000080",
  2884 => x"26089180",
  2885 => x"1d000400",
  2886 => x"1c000000",
  2887 => x"25000000",
  2888 => x"1a000c00",
  2889 => x"1b000000",
  2890 => x"24000000",
  2891 => x"12000000",
  2892 => x"2e000001",
  2893 => x"2d000300",
  2894 => x"23000000",
  2895 => x"36000000",
  2896 => x"21000b00",
  2897 => x"2b000000",
  2898 => x"2c000000",
  2899 => x"22000000",
  2900 => x"3d000000",
  2901 => x"35006c00",
  2902 => x"34000000",
  2903 => x"3e000000",
  2904 => x"32007500",
  2905 => x"33000000",
  2906 => x"3c000000",
  2907 => x"2a006b00",
  2908 => x"46000000",
  2909 => x"43000100",
  2910 => x"3b007300",
  2911 => x"45006900",
  2912 => x"3a000900",
  2913 => x"42007000",
  2914 => x"44007200",
  2915 => x"31007400",
  2916 => x"55000000",
  2917 => x"4d000000",
  2918 => x"4b007c00",
  2919 => x"7b007a00",
  2920 => x"49000000",
  2921 => x"4c007100",
  2922 => x"54008400",
  2923 => x"41007700",
  2924 => x"61000000",
  2925 => x"5b000000",
  2926 => x"52007c00",
  2927 => x"f1000000",
  2928 => x"59000000",
  2929 => x"0e000002",
  2930 => x"5d005d00",
  2931 => x"4a000000",
  2932 => x"16007900",
  2933 => x"76000500",
  2934 => x"0d000700",
  2935 => x"1e000d00",
  2936 => x"29000600",
  2937 => x"14000000",
  2938 => x"15000004",
  2939 => x"00000000",
  2940 => x"00000040",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
