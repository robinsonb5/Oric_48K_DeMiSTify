
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"7f",x"7f",x"30",x"18"),
     1 => (x"36",x"63",x"41",x"00"),
     2 => (x"63",x"36",x"1c",x"1c"),
     3 => (x"06",x"03",x"01",x"41"),
     4 => (x"03",x"06",x"7c",x"7c"),
     5 => (x"59",x"71",x"61",x"01"),
     6 => (x"41",x"43",x"47",x"4d"),
     7 => (x"7f",x"00",x"00",x"00"),
     8 => (x"00",x"41",x"41",x"7f"),
     9 => (x"06",x"03",x"01",x"00"),
    10 => (x"60",x"30",x"18",x"0c"),
    11 => (x"41",x"00",x"00",x"40"),
    12 => (x"00",x"7f",x"7f",x"41"),
    13 => (x"06",x"0c",x"08",x"00"),
    14 => (x"08",x"0c",x"06",x"03"),
    15 => (x"80",x"80",x"80",x"00"),
    16 => (x"80",x"80",x"80",x"80"),
    17 => (x"00",x"00",x"00",x"00"),
    18 => (x"00",x"04",x"07",x"03"),
    19 => (x"74",x"20",x"00",x"00"),
    20 => (x"78",x"7c",x"54",x"54"),
    21 => (x"7f",x"7f",x"00",x"00"),
    22 => (x"38",x"7c",x"44",x"44"),
    23 => (x"7c",x"38",x"00",x"00"),
    24 => (x"00",x"44",x"44",x"44"),
    25 => (x"7c",x"38",x"00",x"00"),
    26 => (x"7f",x"7f",x"44",x"44"),
    27 => (x"7c",x"38",x"00",x"00"),
    28 => (x"18",x"5c",x"54",x"54"),
    29 => (x"7e",x"04",x"00",x"00"),
    30 => (x"00",x"05",x"05",x"7f"),
    31 => (x"bc",x"18",x"00",x"00"),
    32 => (x"7c",x"fc",x"a4",x"a4"),
    33 => (x"7f",x"7f",x"00",x"00"),
    34 => (x"78",x"7c",x"04",x"04"),
    35 => (x"00",x"00",x"00",x"00"),
    36 => (x"00",x"40",x"7d",x"3d"),
    37 => (x"80",x"80",x"00",x"00"),
    38 => (x"00",x"7d",x"fd",x"80"),
    39 => (x"7f",x"7f",x"00",x"00"),
    40 => (x"44",x"6c",x"38",x"10"),
    41 => (x"00",x"00",x"00",x"00"),
    42 => (x"00",x"40",x"7f",x"3f"),
    43 => (x"0c",x"7c",x"7c",x"00"),
    44 => (x"78",x"7c",x"0c",x"18"),
    45 => (x"7c",x"7c",x"00",x"00"),
    46 => (x"78",x"7c",x"04",x"04"),
    47 => (x"7c",x"38",x"00",x"00"),
    48 => (x"38",x"7c",x"44",x"44"),
    49 => (x"fc",x"fc",x"00",x"00"),
    50 => (x"18",x"3c",x"24",x"24"),
    51 => (x"3c",x"18",x"00",x"00"),
    52 => (x"fc",x"fc",x"24",x"24"),
    53 => (x"7c",x"7c",x"00",x"00"),
    54 => (x"08",x"0c",x"04",x"04"),
    55 => (x"5c",x"48",x"00",x"00"),
    56 => (x"20",x"74",x"54",x"54"),
    57 => (x"3f",x"04",x"00",x"00"),
    58 => (x"00",x"44",x"44",x"7f"),
    59 => (x"7c",x"3c",x"00",x"00"),
    60 => (x"7c",x"7c",x"40",x"40"),
    61 => (x"3c",x"1c",x"00",x"00"),
    62 => (x"1c",x"3c",x"60",x"60"),
    63 => (x"60",x"7c",x"3c",x"00"),
    64 => (x"3c",x"7c",x"60",x"30"),
    65 => (x"38",x"6c",x"44",x"00"),
    66 => (x"44",x"6c",x"38",x"10"),
    67 => (x"bc",x"1c",x"00",x"00"),
    68 => (x"1c",x"3c",x"60",x"e0"),
    69 => (x"64",x"44",x"00",x"00"),
    70 => (x"44",x"4c",x"5c",x"74"),
    71 => (x"08",x"08",x"00",x"00"),
    72 => (x"41",x"41",x"77",x"3e"),
    73 => (x"00",x"00",x"00",x"00"),
    74 => (x"00",x"00",x"7f",x"7f"),
    75 => (x"41",x"41",x"00",x"00"),
    76 => (x"08",x"08",x"3e",x"77"),
    77 => (x"01",x"01",x"02",x"00"),
    78 => (x"01",x"02",x"02",x"03"),
    79 => (x"7f",x"7f",x"7f",x"00"),
    80 => (x"7f",x"7f",x"7f",x"7f"),
    81 => (x"1c",x"08",x"08",x"00"),
    82 => (x"7f",x"3e",x"3e",x"1c"),
    83 => (x"3e",x"7f",x"7f",x"7f"),
    84 => (x"08",x"1c",x"1c",x"3e"),
    85 => (x"18",x"10",x"00",x"08"),
    86 => (x"10",x"18",x"7c",x"7c"),
    87 => (x"30",x"10",x"00",x"00"),
    88 => (x"10",x"30",x"7c",x"7c"),
    89 => (x"60",x"30",x"10",x"00"),
    90 => (x"06",x"1e",x"78",x"60"),
    91 => (x"3c",x"66",x"42",x"00"),
    92 => (x"42",x"66",x"3c",x"18"),
    93 => (x"6a",x"38",x"78",x"00"),
    94 => (x"38",x"6c",x"c6",x"c2"),
    95 => (x"00",x"00",x"60",x"00"),
    96 => (x"60",x"00",x"00",x"60"),
    97 => (x"5b",x"5e",x"0e",x"00"),
    98 => (x"1e",x"0e",x"5d",x"5c"),
    99 => (x"c9",x"c3",x"4c",x"71"),
   100 => (x"c0",x"4d",x"bf",x"e2"),
   101 => (x"74",x"1e",x"c0",x"4b"),
   102 => (x"87",x"c7",x"02",x"ab"),
   103 => (x"c0",x"48",x"a6",x"c4"),
   104 => (x"c4",x"87",x"c5",x"78"),
   105 => (x"78",x"c1",x"48",x"a6"),
   106 => (x"73",x"1e",x"66",x"c4"),
   107 => (x"87",x"df",x"ee",x"49"),
   108 => (x"e0",x"c0",x"86",x"c8"),
   109 => (x"87",x"ef",x"ef",x"49"),
   110 => (x"6a",x"4a",x"a5",x"c4"),
   111 => (x"87",x"f0",x"f0",x"49"),
   112 => (x"cb",x"87",x"c6",x"f1"),
   113 => (x"c8",x"83",x"c1",x"85"),
   114 => (x"ff",x"04",x"ab",x"b7"),
   115 => (x"26",x"26",x"87",x"c7"),
   116 => (x"26",x"4c",x"26",x"4d"),
   117 => (x"1e",x"4f",x"26",x"4b"),
   118 => (x"c9",x"c3",x"4a",x"71"),
   119 => (x"c9",x"c3",x"5a",x"e6"),
   120 => (x"78",x"c7",x"48",x"e6"),
   121 => (x"87",x"dd",x"fe",x"49"),
   122 => (x"73",x"1e",x"4f",x"26"),
   123 => (x"c0",x"4a",x"71",x"1e"),
   124 => (x"d3",x"03",x"aa",x"b7"),
   125 => (x"f8",x"d7",x"c2",x"87"),
   126 => (x"87",x"c4",x"05",x"bf"),
   127 => (x"87",x"c2",x"4b",x"c1"),
   128 => (x"d7",x"c2",x"4b",x"c0"),
   129 => (x"87",x"c4",x"5b",x"fc"),
   130 => (x"5a",x"fc",x"d7",x"c2"),
   131 => (x"bf",x"f8",x"d7",x"c2"),
   132 => (x"c1",x"9a",x"c1",x"4a"),
   133 => (x"ec",x"49",x"a2",x"c0"),
   134 => (x"d7",x"c2",x"87",x"e8"),
   135 => (x"c2",x"49",x"bf",x"e0"),
   136 => (x"b1",x"bf",x"f8",x"d7"),
   137 => (x"78",x"71",x"48",x"fc"),
   138 => (x"1e",x"87",x"e8",x"fe"),
   139 => (x"66",x"c4",x"4a",x"71"),
   140 => (x"e9",x"49",x"72",x"1e"),
   141 => (x"26",x"26",x"87",x"f6"),
   142 => (x"d7",x"c2",x"1e",x"4f"),
   143 => (x"c0",x"49",x"bf",x"f8"),
   144 => (x"c3",x"87",x"d7",x"e9"),
   145 => (x"e8",x"48",x"da",x"c9"),
   146 => (x"c9",x"c3",x"78",x"bf"),
   147 => (x"bf",x"ec",x"48",x"d6"),
   148 => (x"da",x"c9",x"c3",x"78"),
   149 => (x"c3",x"49",x"4a",x"bf"),
   150 => (x"b7",x"c8",x"99",x"ff"),
   151 => (x"71",x"48",x"72",x"2a"),
   152 => (x"e2",x"c9",x"c3",x"b0"),
   153 => (x"0e",x"4f",x"26",x"58"),
   154 => (x"5d",x"5c",x"5b",x"5e"),
   155 => (x"ff",x"4b",x"71",x"0e"),
   156 => (x"c9",x"c3",x"87",x"c7"),
   157 => (x"50",x"c0",x"48",x"d5"),
   158 => (x"f5",x"e5",x"49",x"73"),
   159 => (x"4c",x"49",x"70",x"87"),
   160 => (x"ee",x"cb",x"9c",x"c2"),
   161 => (x"87",x"f8",x"cd",x"49"),
   162 => (x"c3",x"4d",x"49",x"70"),
   163 => (x"bf",x"97",x"d5",x"c9"),
   164 => (x"87",x"e2",x"c1",x"05"),
   165 => (x"c3",x"49",x"66",x"d0"),
   166 => (x"99",x"bf",x"de",x"c9"),
   167 => (x"d4",x"87",x"d6",x"05"),
   168 => (x"c9",x"c3",x"49",x"66"),
   169 => (x"05",x"99",x"bf",x"d6"),
   170 => (x"49",x"73",x"87",x"cb"),
   171 => (x"70",x"87",x"c3",x"e5"),
   172 => (x"c1",x"c1",x"02",x"98"),
   173 => (x"fd",x"4c",x"c1",x"87"),
   174 => (x"49",x"75",x"87",x"ff"),
   175 => (x"70",x"87",x"cd",x"cd"),
   176 => (x"87",x"c6",x"02",x"98"),
   177 => (x"48",x"d5",x"c9",x"c3"),
   178 => (x"c9",x"c3",x"50",x"c1"),
   179 => (x"05",x"bf",x"97",x"d5"),
   180 => (x"c3",x"87",x"e3",x"c0"),
   181 => (x"49",x"bf",x"de",x"c9"),
   182 => (x"05",x"99",x"66",x"d0"),
   183 => (x"c3",x"87",x"d6",x"ff"),
   184 => (x"49",x"bf",x"d6",x"c9"),
   185 => (x"05",x"99",x"66",x"d4"),
   186 => (x"73",x"87",x"ca",x"ff"),
   187 => (x"87",x"c2",x"e4",x"49"),
   188 => (x"fe",x"05",x"98",x"70"),
   189 => (x"48",x"74",x"87",x"ff"),
   190 => (x"0e",x"87",x"d4",x"fb"),
   191 => (x"5d",x"5c",x"5b",x"5e"),
   192 => (x"c0",x"86",x"f8",x"0e"),
   193 => (x"bf",x"ec",x"4c",x"4d"),
   194 => (x"48",x"a6",x"c4",x"7e"),
   195 => (x"bf",x"e2",x"c9",x"c3"),
   196 => (x"1e",x"1e",x"c0",x"78"),
   197 => (x"fd",x"49",x"f7",x"c1"),
   198 => (x"86",x"c8",x"87",x"cd"),
   199 => (x"c0",x"02",x"98",x"70"),
   200 => (x"d7",x"c2",x"87",x"f3"),
   201 => (x"c4",x"05",x"bf",x"e0"),
   202 => (x"c2",x"7e",x"c1",x"87"),
   203 => (x"c2",x"7e",x"c0",x"87"),
   204 => (x"6e",x"48",x"e0",x"d7"),
   205 => (x"1e",x"fc",x"ca",x"78"),
   206 => (x"c9",x"02",x"66",x"c4"),
   207 => (x"48",x"a6",x"c4",x"87"),
   208 => (x"78",x"f7",x"d5",x"c2"),
   209 => (x"a6",x"c4",x"87",x"c7"),
   210 => (x"c2",x"d6",x"c2",x"48"),
   211 => (x"49",x"66",x"c4",x"78"),
   212 => (x"c4",x"87",x"fb",x"c8"),
   213 => (x"c0",x"1e",x"c1",x"86"),
   214 => (x"fc",x"49",x"c7",x"1e"),
   215 => (x"86",x"c8",x"87",x"c9"),
   216 => (x"cd",x"02",x"98",x"70"),
   217 => (x"fa",x"49",x"ff",x"87"),
   218 => (x"da",x"c1",x"87",x"c0"),
   219 => (x"87",x"c2",x"e2",x"49"),
   220 => (x"c9",x"c3",x"4d",x"c1"),
   221 => (x"02",x"bf",x"97",x"d5"),
   222 => (x"f4",x"d6",x"87",x"c3"),
   223 => (x"da",x"c9",x"c3",x"87"),
   224 => (x"d7",x"c2",x"4b",x"bf"),
   225 => (x"c1",x"05",x"bf",x"f8"),
   226 => (x"d7",x"c2",x"87",x"e1"),
   227 => (x"c0",x"02",x"bf",x"e0"),
   228 => (x"a6",x"c4",x"87",x"f0"),
   229 => (x"c0",x"c0",x"c8",x"48"),
   230 => (x"e4",x"d7",x"c2",x"78"),
   231 => (x"bf",x"97",x"6e",x"7e"),
   232 => (x"c1",x"48",x"6e",x"49"),
   233 => (x"71",x"7e",x"70",x"80"),
   234 => (x"70",x"87",x"c7",x"e1"),
   235 => (x"87",x"c3",x"02",x"98"),
   236 => (x"c4",x"b3",x"66",x"c4"),
   237 => (x"b7",x"c1",x"48",x"66"),
   238 => (x"58",x"a6",x"c8",x"28"),
   239 => (x"ff",x"05",x"98",x"70"),
   240 => (x"fd",x"c3",x"87",x"db"),
   241 => (x"87",x"ea",x"e0",x"49"),
   242 => (x"e0",x"49",x"fa",x"c3"),
   243 => (x"49",x"73",x"87",x"e4"),
   244 => (x"71",x"99",x"ff",x"c3"),
   245 => (x"f9",x"49",x"c0",x"1e"),
   246 => (x"49",x"73",x"87",x"d1"),
   247 => (x"71",x"29",x"b7",x"c8"),
   248 => (x"f9",x"49",x"c1",x"1e"),
   249 => (x"86",x"c8",x"87",x"c5"),
   250 => (x"c3",x"87",x"c7",x"c6"),
   251 => (x"4b",x"bf",x"de",x"c9"),
   252 => (x"87",x"df",x"02",x"9b"),
   253 => (x"bf",x"f4",x"d7",x"c2"),
   254 => (x"87",x"d0",x"c8",x"49"),
   255 => (x"c0",x"05",x"98",x"70"),
   256 => (x"4b",x"c0",x"87",x"c4"),
   257 => (x"e0",x"c2",x"87",x"d3"),
   258 => (x"87",x"f4",x"c7",x"49"),
   259 => (x"58",x"f8",x"d7",x"c2"),
   260 => (x"c2",x"87",x"c6",x"c0"),
   261 => (x"c0",x"48",x"f4",x"d7"),
   262 => (x"c2",x"49",x"73",x"78"),
   263 => (x"cf",x"c0",x"05",x"99"),
   264 => (x"49",x"eb",x"c3",x"87"),
   265 => (x"87",x"ca",x"df",x"ff"),
   266 => (x"99",x"c2",x"49",x"70"),
   267 => (x"87",x"c2",x"c0",x"02"),
   268 => (x"49",x"73",x"4c",x"fb"),
   269 => (x"c0",x"05",x"99",x"c1"),
   270 => (x"f4",x"c3",x"87",x"cf"),
   271 => (x"f1",x"de",x"ff",x"49"),
   272 => (x"c2",x"49",x"70",x"87"),
   273 => (x"c2",x"c0",x"02",x"99"),
   274 => (x"73",x"4c",x"fa",x"87"),
   275 => (x"05",x"99",x"c8",x"49"),
   276 => (x"c3",x"87",x"cf",x"c0"),
   277 => (x"de",x"ff",x"49",x"f5"),
   278 => (x"49",x"70",x"87",x"d8"),
   279 => (x"c0",x"02",x"99",x"c2"),
   280 => (x"c9",x"c3",x"87",x"d6"),
   281 => (x"c0",x"02",x"bf",x"e6"),
   282 => (x"c1",x"48",x"87",x"ca"),
   283 => (x"ea",x"c9",x"c3",x"88"),
   284 => (x"87",x"c2",x"c0",x"58"),
   285 => (x"4d",x"c1",x"4c",x"ff"),
   286 => (x"99",x"c4",x"49",x"73"),
   287 => (x"87",x"cf",x"c0",x"05"),
   288 => (x"ff",x"49",x"f2",x"c3"),
   289 => (x"70",x"87",x"eb",x"dd"),
   290 => (x"02",x"99",x"c2",x"49"),
   291 => (x"c3",x"87",x"dc",x"c0"),
   292 => (x"7e",x"bf",x"e6",x"c9"),
   293 => (x"a8",x"b7",x"c7",x"48"),
   294 => (x"87",x"cb",x"c0",x"03"),
   295 => (x"80",x"c1",x"48",x"6e"),
   296 => (x"58",x"ea",x"c9",x"c3"),
   297 => (x"fe",x"87",x"c2",x"c0"),
   298 => (x"c3",x"4d",x"c1",x"4c"),
   299 => (x"dd",x"ff",x"49",x"fd"),
   300 => (x"49",x"70",x"87",x"c0"),
   301 => (x"c0",x"02",x"99",x"c2"),
   302 => (x"c9",x"c3",x"87",x"d5"),
   303 => (x"c0",x"02",x"bf",x"e6"),
   304 => (x"c9",x"c3",x"87",x"c9"),
   305 => (x"78",x"c0",x"48",x"e6"),
   306 => (x"fd",x"87",x"c2",x"c0"),
   307 => (x"c3",x"4d",x"c1",x"4c"),
   308 => (x"dc",x"ff",x"49",x"fa"),
   309 => (x"49",x"70",x"87",x"dc"),
   310 => (x"c0",x"02",x"99",x"c2"),
   311 => (x"c9",x"c3",x"87",x"d9"),
   312 => (x"c7",x"48",x"bf",x"e6"),
   313 => (x"c0",x"03",x"a8",x"b7"),
   314 => (x"c9",x"c3",x"87",x"c9"),
   315 => (x"78",x"c7",x"48",x"e6"),
   316 => (x"fc",x"87",x"c2",x"c0"),
   317 => (x"c0",x"4d",x"c1",x"4c"),
   318 => (x"c0",x"03",x"ac",x"b7"),
   319 => (x"66",x"c4",x"87",x"d5"),
   320 => (x"80",x"d8",x"c1",x"48"),
   321 => (x"bf",x"6e",x"7e",x"70"),
   322 => (x"87",x"c7",x"c0",x"02"),
   323 => (x"74",x"4b",x"bf",x"6e"),
   324 => (x"c0",x"0f",x"73",x"49"),
   325 => (x"1e",x"f0",x"c3",x"1e"),
   326 => (x"f5",x"49",x"da",x"c1"),
   327 => (x"86",x"c8",x"87",x"c9"),
   328 => (x"c0",x"02",x"98",x"70"),
   329 => (x"c9",x"c3",x"87",x"d9"),
   330 => (x"6e",x"7e",x"bf",x"e6"),
   331 => (x"c4",x"91",x"cb",x"49"),
   332 => (x"82",x"71",x"4a",x"66"),
   333 => (x"c6",x"c0",x"02",x"6a"),
   334 => (x"6e",x"4b",x"6a",x"87"),
   335 => (x"75",x"0f",x"73",x"49"),
   336 => (x"c8",x"c0",x"02",x"9d"),
   337 => (x"e6",x"c9",x"c3",x"87"),
   338 => (x"f8",x"f0",x"49",x"bf"),
   339 => (x"fc",x"d7",x"c2",x"87"),
   340 => (x"dd",x"c0",x"02",x"bf"),
   341 => (x"f3",x"c2",x"49",x"87"),
   342 => (x"02",x"98",x"70",x"87"),
   343 => (x"c3",x"87",x"d3",x"c0"),
   344 => (x"49",x"bf",x"e6",x"c9"),
   345 => (x"c0",x"87",x"de",x"f0"),
   346 => (x"87",x"fe",x"f1",x"49"),
   347 => (x"48",x"fc",x"d7",x"c2"),
   348 => (x"8e",x"f8",x"78",x"c0"),
   349 => (x"4a",x"87",x"d8",x"f1"),
   350 => (x"65",x"6b",x"79",x"6f"),
   351 => (x"6f",x"20",x"73",x"79"),
   352 => (x"6f",x"4a",x"00",x"6e"),
   353 => (x"79",x"65",x"6b",x"79"),
   354 => (x"66",x"6f",x"20",x"73"),
   355 => (x"5e",x"0e",x"00",x"66"),
   356 => (x"0e",x"5d",x"5c",x"5b"),
   357 => (x"c3",x"4c",x"71",x"1e"),
   358 => (x"49",x"bf",x"e2",x"c9"),
   359 => (x"4d",x"a1",x"cd",x"c1"),
   360 => (x"69",x"81",x"d1",x"c1"),
   361 => (x"02",x"9c",x"74",x"7e"),
   362 => (x"a5",x"c4",x"87",x"cf"),
   363 => (x"c3",x"7b",x"74",x"4b"),
   364 => (x"49",x"bf",x"e2",x"c9"),
   365 => (x"6e",x"87",x"e0",x"f0"),
   366 => (x"05",x"9c",x"74",x"7b"),
   367 => (x"4b",x"c0",x"87",x"c4"),
   368 => (x"4b",x"c1",x"87",x"c2"),
   369 => (x"e1",x"f0",x"49",x"73"),
   370 => (x"02",x"66",x"d4",x"87"),
   371 => (x"c0",x"49",x"87",x"c8"),
   372 => (x"4a",x"70",x"87",x"ee"),
   373 => (x"4a",x"c0",x"87",x"c2"),
   374 => (x"5a",x"c0",x"d8",x"c2"),
   375 => (x"87",x"ef",x"ef",x"26"),
   376 => (x"00",x"00",x"00",x"00"),
   377 => (x"14",x"11",x"12",x"58"),
   378 => (x"23",x"1c",x"1b",x"1d"),
   379 => (x"94",x"91",x"59",x"5a"),
   380 => (x"f4",x"eb",x"f2",x"f5"),
   381 => (x"00",x"00",x"00",x"00"),
   382 => (x"00",x"00",x"00",x"00"),
   383 => (x"00",x"00",x"00",x"00"),
   384 => (x"ff",x"4a",x"71",x"1e"),
   385 => (x"72",x"49",x"bf",x"c8"),
   386 => (x"4f",x"26",x"48",x"a1"),
   387 => (x"bf",x"c8",x"ff",x"1e"),
   388 => (x"c0",x"c0",x"fe",x"89"),
   389 => (x"a9",x"c0",x"c0",x"c0"),
   390 => (x"c0",x"87",x"c4",x"01"),
   391 => (x"c1",x"87",x"c2",x"4a"),
   392 => (x"26",x"48",x"72",x"4a"),
   393 => (x"5b",x"5e",x"0e",x"4f"),
   394 => (x"71",x"0e",x"5d",x"5c"),
   395 => (x"4c",x"d4",x"ff",x"4b"),
   396 => (x"c0",x"48",x"66",x"d0"),
   397 => (x"ff",x"49",x"d6",x"78"),
   398 => (x"c3",x"87",x"f7",x"d8"),
   399 => (x"49",x"6c",x"7c",x"ff"),
   400 => (x"71",x"99",x"ff",x"c3"),
   401 => (x"f0",x"c3",x"49",x"4d"),
   402 => (x"a9",x"e0",x"c1",x"99"),
   403 => (x"c3",x"87",x"cb",x"05"),
   404 => (x"48",x"6c",x"7c",x"ff"),
   405 => (x"66",x"d0",x"98",x"c3"),
   406 => (x"ff",x"c3",x"78",x"08"),
   407 => (x"49",x"4a",x"6c",x"7c"),
   408 => (x"ff",x"c3",x"31",x"c8"),
   409 => (x"71",x"4a",x"6c",x"7c"),
   410 => (x"c8",x"49",x"72",x"b2"),
   411 => (x"7c",x"ff",x"c3",x"31"),
   412 => (x"b2",x"71",x"4a",x"6c"),
   413 => (x"31",x"c8",x"49",x"72"),
   414 => (x"6c",x"7c",x"ff",x"c3"),
   415 => (x"ff",x"b2",x"71",x"4a"),
   416 => (x"e0",x"c0",x"48",x"d0"),
   417 => (x"02",x"9b",x"73",x"78"),
   418 => (x"7b",x"72",x"87",x"c2"),
   419 => (x"4d",x"26",x"48",x"75"),
   420 => (x"4b",x"26",x"4c",x"26"),
   421 => (x"26",x"1e",x"4f",x"26"),
   422 => (x"5b",x"5e",x"0e",x"4f"),
   423 => (x"86",x"f8",x"0e",x"5c"),
   424 => (x"a6",x"c8",x"1e",x"76"),
   425 => (x"87",x"fd",x"fd",x"49"),
   426 => (x"4b",x"70",x"86",x"c4"),
   427 => (x"a8",x"c2",x"48",x"6e"),
   428 => (x"87",x"ca",x"c3",x"03"),
   429 => (x"f0",x"c3",x"4a",x"73"),
   430 => (x"aa",x"d0",x"c1",x"9a"),
   431 => (x"c1",x"87",x"c7",x"02"),
   432 => (x"c2",x"05",x"aa",x"e0"),
   433 => (x"49",x"73",x"87",x"f8"),
   434 => (x"c3",x"02",x"99",x"c8"),
   435 => (x"87",x"c6",x"ff",x"87"),
   436 => (x"9c",x"c3",x"4c",x"73"),
   437 => (x"c1",x"05",x"ac",x"c2"),
   438 => (x"66",x"c4",x"87",x"cf"),
   439 => (x"71",x"31",x"c9",x"49"),
   440 => (x"4a",x"66",x"c4",x"1e"),
   441 => (x"c3",x"92",x"c8",x"c1"),
   442 => (x"72",x"49",x"ea",x"c9"),
   443 => (x"de",x"d0",x"fe",x"81"),
   444 => (x"49",x"66",x"c4",x"87"),
   445 => (x"49",x"e3",x"c0",x"1e"),
   446 => (x"87",x"db",x"d6",x"ff"),
   447 => (x"d5",x"ff",x"49",x"d8"),
   448 => (x"c0",x"c8",x"87",x"f0"),
   449 => (x"da",x"f8",x"c2",x"1e"),
   450 => (x"f3",x"e8",x"fd",x"49"),
   451 => (x"48",x"d0",x"ff",x"87"),
   452 => (x"c2",x"78",x"e0",x"c0"),
   453 => (x"d0",x"1e",x"da",x"f8"),
   454 => (x"c8",x"c1",x"4a",x"66"),
   455 => (x"ea",x"c9",x"c3",x"92"),
   456 => (x"fe",x"81",x"72",x"49"),
   457 => (x"d0",x"87",x"e6",x"cb"),
   458 => (x"05",x"ac",x"c1",x"86"),
   459 => (x"c4",x"87",x"cf",x"c1"),
   460 => (x"31",x"c9",x"49",x"66"),
   461 => (x"66",x"c4",x"1e",x"71"),
   462 => (x"92",x"c8",x"c1",x"4a"),
   463 => (x"49",x"ea",x"c9",x"c3"),
   464 => (x"cf",x"fe",x"81",x"72"),
   465 => (x"f8",x"c2",x"87",x"c9"),
   466 => (x"66",x"c8",x"1e",x"da"),
   467 => (x"92",x"c8",x"c1",x"4a"),
   468 => (x"49",x"ea",x"c9",x"c3"),
   469 => (x"c9",x"fe",x"81",x"72"),
   470 => (x"66",x"c8",x"87",x"f0"),
   471 => (x"e3",x"c0",x"1e",x"49"),
   472 => (x"f2",x"d4",x"ff",x"49"),
   473 => (x"ff",x"49",x"d7",x"87"),
   474 => (x"c8",x"87",x"c7",x"d4"),
   475 => (x"f8",x"c2",x"1e",x"c0"),
   476 => (x"e6",x"fd",x"49",x"da"),
   477 => (x"86",x"d0",x"87",x"f4"),
   478 => (x"c0",x"48",x"d0",x"ff"),
   479 => (x"8e",x"f8",x"78",x"e0"),
   480 => (x"0e",x"87",x"cd",x"fc"),
   481 => (x"5d",x"5c",x"5b",x"5e"),
   482 => (x"4d",x"71",x"1e",x"0e"),
   483 => (x"d4",x"4c",x"d4",x"ff"),
   484 => (x"c3",x"48",x"7e",x"66"),
   485 => (x"c5",x"06",x"a8",x"b7"),
   486 => (x"c1",x"48",x"c0",x"87"),
   487 => (x"49",x"75",x"87",x"e3"),
   488 => (x"87",x"d2",x"df",x"fe"),
   489 => (x"66",x"c4",x"1e",x"75"),
   490 => (x"93",x"c8",x"c1",x"4b"),
   491 => (x"83",x"ea",x"c9",x"c3"),
   492 => (x"c3",x"fe",x"49",x"73"),
   493 => (x"83",x"c8",x"87",x"fe"),
   494 => (x"d0",x"ff",x"4b",x"6b"),
   495 => (x"78",x"e1",x"c8",x"48"),
   496 => (x"49",x"73",x"7c",x"dd"),
   497 => (x"71",x"99",x"ff",x"c3"),
   498 => (x"c8",x"49",x"73",x"7c"),
   499 => (x"ff",x"c3",x"29",x"b7"),
   500 => (x"73",x"7c",x"71",x"99"),
   501 => (x"29",x"b7",x"d0",x"49"),
   502 => (x"71",x"99",x"ff",x"c3"),
   503 => (x"d8",x"49",x"73",x"7c"),
   504 => (x"7c",x"71",x"29",x"b7"),
   505 => (x"7c",x"7c",x"7c",x"c0"),
   506 => (x"7c",x"7c",x"7c",x"7c"),
   507 => (x"7c",x"7c",x"7c",x"7c"),
   508 => (x"78",x"e0",x"c0",x"7c"),
   509 => (x"dc",x"1e",x"66",x"c4"),
   510 => (x"da",x"d2",x"ff",x"49"),
   511 => (x"73",x"86",x"c8",x"87"),
   512 => (x"c9",x"fa",x"26",x"48"),
   513 => (x"5b",x"5e",x"0e",x"87"),
   514 => (x"1e",x"0e",x"5d",x"5c"),
   515 => (x"d4",x"ff",x"7e",x"71"),
   516 => (x"c3",x"1e",x"6e",x"4b"),
   517 => (x"fe",x"49",x"fa",x"cb"),
   518 => (x"c4",x"87",x"d9",x"c2"),
   519 => (x"9d",x"4d",x"70",x"86"),
   520 => (x"87",x"c3",x"c3",x"02"),
   521 => (x"bf",x"c2",x"cc",x"c3"),
   522 => (x"fe",x"49",x"6e",x"4c"),
   523 => (x"ff",x"87",x"c7",x"dd"),
   524 => (x"c5",x"c8",x"48",x"d0"),
   525 => (x"7b",x"d6",x"c1",x"78"),
   526 => (x"7b",x"15",x"4a",x"c0"),
   527 => (x"e0",x"c0",x"82",x"c1"),
   528 => (x"f5",x"04",x"aa",x"b7"),
   529 => (x"48",x"d0",x"ff",x"87"),
   530 => (x"c5",x"c8",x"78",x"c4"),
   531 => (x"7b",x"d3",x"c1",x"78"),
   532 => (x"78",x"c4",x"7b",x"c1"),
   533 => (x"c1",x"02",x"9c",x"74"),
   534 => (x"f8",x"c2",x"87",x"fc"),
   535 => (x"c0",x"c8",x"7e",x"da"),
   536 => (x"b7",x"c0",x"8c",x"4d"),
   537 => (x"87",x"c6",x"03",x"ac"),
   538 => (x"4d",x"a4",x"c0",x"c8"),
   539 => (x"c5",x"c3",x"4c",x"c0"),
   540 => (x"49",x"bf",x"97",x"cb"),
   541 => (x"d2",x"02",x"99",x"d0"),
   542 => (x"c3",x"1e",x"c0",x"87"),
   543 => (x"fe",x"49",x"fa",x"cb"),
   544 => (x"c4",x"87",x"c7",x"c5"),
   545 => (x"4a",x"49",x"70",x"86"),
   546 => (x"c2",x"87",x"ef",x"c0"),
   547 => (x"c3",x"1e",x"da",x"f8"),
   548 => (x"fe",x"49",x"fa",x"cb"),
   549 => (x"c4",x"87",x"f3",x"c4"),
   550 => (x"4a",x"49",x"70",x"86"),
   551 => (x"c8",x"48",x"d0",x"ff"),
   552 => (x"d4",x"c1",x"78",x"c5"),
   553 => (x"bf",x"97",x"6e",x"7b"),
   554 => (x"c1",x"48",x"6e",x"7b"),
   555 => (x"c1",x"7e",x"70",x"80"),
   556 => (x"f0",x"ff",x"05",x"8d"),
   557 => (x"48",x"d0",x"ff",x"87"),
   558 => (x"9a",x"72",x"78",x"c4"),
   559 => (x"c0",x"87",x"c5",x"05"),
   560 => (x"87",x"e5",x"c0",x"48"),
   561 => (x"cb",x"c3",x"1e",x"c1"),
   562 => (x"c2",x"fe",x"49",x"fa"),
   563 => (x"86",x"c4",x"87",x"db"),
   564 => (x"fe",x"05",x"9c",x"74"),
   565 => (x"d0",x"ff",x"87",x"c4"),
   566 => (x"78",x"c5",x"c8",x"48"),
   567 => (x"c0",x"7b",x"d3",x"c1"),
   568 => (x"c1",x"78",x"c4",x"7b"),
   569 => (x"c0",x"87",x"c2",x"48"),
   570 => (x"4d",x"26",x"26",x"48"),
   571 => (x"4b",x"26",x"4c",x"26"),
   572 => (x"5e",x"0e",x"4f",x"26"),
   573 => (x"71",x"0e",x"5c",x"5b"),
   574 => (x"02",x"66",x"cc",x"4b"),
   575 => (x"c0",x"4c",x"87",x"d8"),
   576 => (x"d8",x"02",x"8c",x"f0"),
   577 => (x"c1",x"4a",x"74",x"87"),
   578 => (x"87",x"d1",x"02",x"8a"),
   579 => (x"87",x"cd",x"02",x"8a"),
   580 => (x"87",x"c9",x"02",x"8a"),
   581 => (x"49",x"73",x"87",x"d7"),
   582 => (x"d0",x"87",x"ea",x"fb"),
   583 => (x"c0",x"1e",x"74",x"87"),
   584 => (x"87",x"df",x"f9",x"49"),
   585 => (x"49",x"73",x"1e",x"74"),
   586 => (x"c8",x"87",x"d8",x"f9"),
   587 => (x"87",x"fc",x"fe",x"86"),
   588 => (x"e5",x"c2",x"1e",x"00"),
   589 => (x"c1",x"49",x"bf",x"da"),
   590 => (x"de",x"e5",x"c2",x"b9"),
   591 => (x"48",x"d4",x"ff",x"59"),
   592 => (x"ff",x"78",x"ff",x"c3"),
   593 => (x"e1",x"c8",x"48",x"d0"),
   594 => (x"48",x"d4",x"ff",x"78"),
   595 => (x"31",x"c4",x"78",x"c1"),
   596 => (x"d0",x"ff",x"78",x"71"),
   597 => (x"78",x"e0",x"c0",x"48"),
   598 => (x"00",x"00",x"4f",x"26"),
   599 => (x"ff",x"1e",x"00",x"00"),
   600 => (x"c4",x"87",x"dd",x"c1"),
   601 => (x"c0",x"c2",x"49",x"66"),
   602 => (x"87",x"cd",x"02",x"99"),
   603 => (x"c3",x"1e",x"e0",x"c3"),
   604 => (x"ff",x"49",x"f7",x"c8"),
   605 => (x"c4",x"87",x"ec",x"c2"),
   606 => (x"49",x"66",x"c4",x"86"),
   607 => (x"02",x"99",x"c0",x"c4"),
   608 => (x"f0",x"c3",x"87",x"cd"),
   609 => (x"f7",x"c8",x"c3",x"1e"),
   610 => (x"d6",x"c2",x"ff",x"49"),
   611 => (x"c4",x"86",x"c4",x"87"),
   612 => (x"ff",x"c1",x"49",x"66"),
   613 => (x"c3",x"1e",x"71",x"99"),
   614 => (x"ff",x"49",x"f7",x"c8"),
   615 => (x"ff",x"87",x"c4",x"c2"),
   616 => (x"26",x"87",x"d5",x"c0"),
   617 => (x"5e",x"0e",x"4f",x"26"),
   618 => (x"0e",x"5d",x"5c",x"5b"),
   619 => (x"c0",x"86",x"d8",x"ff"),
   620 => (x"c6",x"cd",x"c3",x"7e"),
   621 => (x"81",x"c2",x"49",x"bf"),
   622 => (x"1e",x"72",x"1e",x"71"),
   623 => (x"dc",x"fd",x"4a",x"c6"),
   624 => (x"48",x"71",x"87",x"f7"),
   625 => (x"49",x"26",x"4a",x"26"),
   626 => (x"c3",x"58",x"a6",x"c8"),
   627 => (x"49",x"bf",x"c6",x"cd"),
   628 => (x"1e",x"71",x"81",x"c4"),
   629 => (x"4a",x"c6",x"1e",x"72"),
   630 => (x"87",x"dd",x"dc",x"fd"),
   631 => (x"4a",x"26",x"48",x"71"),
   632 => (x"a6",x"cc",x"49",x"26"),
   633 => (x"f7",x"f1",x"c2",x"58"),
   634 => (x"df",x"f0",x"49",x"bf"),
   635 => (x"02",x"98",x"70",x"87"),
   636 => (x"c0",x"87",x"f9",x"c9"),
   637 => (x"c7",x"f0",x"49",x"e0"),
   638 => (x"c2",x"49",x"70",x"87"),
   639 => (x"c0",x"59",x"fb",x"f1"),
   640 => (x"c4",x"49",x"74",x"4c"),
   641 => (x"81",x"d0",x"fe",x"91"),
   642 => (x"49",x"74",x"4a",x"69"),
   643 => (x"bf",x"c6",x"cd",x"c3"),
   644 => (x"c3",x"91",x"c4",x"81"),
   645 => (x"72",x"81",x"d2",x"cd"),
   646 => (x"d2",x"02",x"9a",x"79"),
   647 => (x"c1",x"49",x"72",x"87"),
   648 => (x"6e",x"9a",x"71",x"89"),
   649 => (x"70",x"80",x"c1",x"48"),
   650 => (x"05",x"9a",x"72",x"7e"),
   651 => (x"c1",x"87",x"ee",x"ff"),
   652 => (x"ac",x"b7",x"c2",x"84"),
   653 => (x"87",x"c9",x"ff",x"04"),
   654 => (x"fc",x"c0",x"48",x"6e"),
   655 => (x"c8",x"04",x"a8",x"b7"),
   656 => (x"4c",x"c0",x"87",x"ea"),
   657 => (x"66",x"c4",x"4a",x"74"),
   658 => (x"c3",x"92",x"c4",x"82"),
   659 => (x"74",x"82",x"d2",x"cd"),
   660 => (x"81",x"66",x"c8",x"49"),
   661 => (x"cd",x"c3",x"91",x"c4"),
   662 => (x"4a",x"6a",x"81",x"d2"),
   663 => (x"b9",x"72",x"49",x"69"),
   664 => (x"cd",x"c3",x"4b",x"74"),
   665 => (x"c4",x"83",x"bf",x"c6"),
   666 => (x"d2",x"cd",x"c3",x"93"),
   667 => (x"72",x"ba",x"6b",x"83"),
   668 => (x"d4",x"98",x"71",x"48"),
   669 => (x"49",x"74",x"58",x"a6"),
   670 => (x"bf",x"c6",x"cd",x"c3"),
   671 => (x"c3",x"91",x"c4",x"81"),
   672 => (x"69",x"81",x"d2",x"cd"),
   673 => (x"48",x"a6",x"d4",x"7e"),
   674 => (x"a6",x"d0",x"78",x"c0"),
   675 => (x"4c",x"ff",x"c3",x"5c"),
   676 => (x"df",x"49",x"66",x"d0"),
   677 => (x"e2",x"c6",x"02",x"29"),
   678 => (x"4a",x"66",x"cc",x"87"),
   679 => (x"d4",x"92",x"e0",x"c0"),
   680 => (x"ff",x"c0",x"82",x"66"),
   681 => (x"70",x"88",x"72",x"48"),
   682 => (x"48",x"a6",x"d8",x"4a"),
   683 => (x"80",x"c4",x"78",x"c0"),
   684 => (x"49",x"6e",x"78",x"c0"),
   685 => (x"e4",x"c0",x"29",x"df"),
   686 => (x"cd",x"c3",x"59",x"a6"),
   687 => (x"78",x"c1",x"48",x"c2"),
   688 => (x"31",x"c3",x"49",x"72"),
   689 => (x"b1",x"72",x"2a",x"b7"),
   690 => (x"c4",x"99",x"ff",x"c0"),
   691 => (x"f3",x"f3",x"c2",x"91"),
   692 => (x"6d",x"85",x"71",x"4d"),
   693 => (x"c0",x"c4",x"49",x"4b"),
   694 => (x"d7",x"02",x"99",x"c0"),
   695 => (x"66",x"e0",x"c0",x"87"),
   696 => (x"87",x"c7",x"c0",x"02"),
   697 => (x"78",x"c0",x"80",x"c8"),
   698 => (x"c3",x"87",x"d0",x"c5"),
   699 => (x"c1",x"48",x"ca",x"cd"),
   700 => (x"87",x"c7",x"c5",x"78"),
   701 => (x"02",x"66",x"e0",x"c0"),
   702 => (x"49",x"73",x"87",x"d8"),
   703 => (x"99",x"c0",x"c0",x"c2"),
   704 => (x"87",x"c3",x"c0",x"02"),
   705 => (x"6d",x"2b",x"b7",x"d0"),
   706 => (x"ff",x"ff",x"fd",x"48"),
   707 => (x"c0",x"7d",x"70",x"98"),
   708 => (x"cd",x"c3",x"87",x"fa"),
   709 => (x"c0",x"02",x"bf",x"ca"),
   710 => (x"48",x"73",x"87",x"f2"),
   711 => (x"c0",x"28",x"b7",x"d0"),
   712 => (x"70",x"58",x"a6",x"e8"),
   713 => (x"e3",x"c0",x"02",x"98"),
   714 => (x"ce",x"cd",x"c3",x"87"),
   715 => (x"e0",x"c0",x"49",x"bf"),
   716 => (x"c0",x"02",x"99",x"c0"),
   717 => (x"49",x"70",x"87",x"ca"),
   718 => (x"99",x"c0",x"e0",x"c0"),
   719 => (x"87",x"cc",x"c0",x"02"),
   720 => (x"c0",x"c2",x"48",x"6d"),
   721 => (x"7d",x"70",x"b0",x"c0"),
   722 => (x"4b",x"66",x"e4",x"c0"),
   723 => (x"c0",x"c8",x"49",x"73"),
   724 => (x"c2",x"02",x"99",x"c0"),
   725 => (x"cd",x"c3",x"87",x"c5"),
   726 => (x"cc",x"4a",x"bf",x"ce"),
   727 => (x"c0",x"02",x"9a",x"c0"),
   728 => (x"c0",x"c4",x"87",x"cf"),
   729 => (x"d7",x"c0",x"02",x"8a"),
   730 => (x"c0",x"02",x"8a",x"87"),
   731 => (x"dc",x"c1",x"87",x"f8"),
   732 => (x"74",x"49",x"73",x"87"),
   733 => (x"c2",x"91",x"c2",x"99"),
   734 => (x"11",x"81",x"e7",x"f3"),
   735 => (x"87",x"db",x"c1",x"4b"),
   736 => (x"99",x"74",x"49",x"73"),
   737 => (x"f3",x"c2",x"91",x"c2"),
   738 => (x"81",x"c1",x"81",x"e7"),
   739 => (x"e0",x"c0",x"4b",x"11"),
   740 => (x"c8",x"c0",x"02",x"66"),
   741 => (x"48",x"a6",x"dc",x"87"),
   742 => (x"fe",x"c0",x"78",x"d2"),
   743 => (x"48",x"a6",x"d8",x"87"),
   744 => (x"c0",x"78",x"d2",x"c4"),
   745 => (x"49",x"73",x"87",x"f5"),
   746 => (x"91",x"c2",x"99",x"74"),
   747 => (x"81",x"e7",x"f3",x"c2"),
   748 => (x"4b",x"11",x"81",x"c1"),
   749 => (x"02",x"66",x"e0",x"c0"),
   750 => (x"dc",x"87",x"c9",x"c0"),
   751 => (x"d9",x"c1",x"48",x"a6"),
   752 => (x"87",x"d7",x"c0",x"78"),
   753 => (x"c5",x"48",x"a6",x"d8"),
   754 => (x"ce",x"c0",x"78",x"d9"),
   755 => (x"74",x"49",x"73",x"87"),
   756 => (x"c2",x"91",x"c2",x"99"),
   757 => (x"c1",x"81",x"e7",x"f3"),
   758 => (x"c0",x"4b",x"11",x"81"),
   759 => (x"c0",x"02",x"66",x"e0"),
   760 => (x"49",x"73",x"87",x"db"),
   761 => (x"fc",x"c7",x"b9",x"ff"),
   762 => (x"48",x"71",x"99",x"c0"),
   763 => (x"bf",x"ce",x"cd",x"c3"),
   764 => (x"d2",x"cd",x"c3",x"98"),
   765 => (x"c4",x"9b",x"74",x"58"),
   766 => (x"d3",x"c0",x"b3",x"c0"),
   767 => (x"c7",x"49",x"73",x"87"),
   768 => (x"71",x"99",x"c0",x"fc"),
   769 => (x"ce",x"cd",x"c3",x"48"),
   770 => (x"cd",x"c3",x"b0",x"bf"),
   771 => (x"9b",x"74",x"58",x"d2"),
   772 => (x"c0",x"02",x"66",x"d8"),
   773 => (x"c3",x"1e",x"87",x"ca"),
   774 => (x"f5",x"49",x"c2",x"cd"),
   775 => (x"86",x"c4",x"87",x"c0"),
   776 => (x"cd",x"c3",x"1e",x"73"),
   777 => (x"f5",x"f4",x"49",x"c2"),
   778 => (x"dc",x"86",x"c4",x"87"),
   779 => (x"ca",x"c0",x"02",x"66"),
   780 => (x"cd",x"c3",x"1e",x"87"),
   781 => (x"e5",x"f4",x"49",x"c2"),
   782 => (x"d0",x"86",x"c4",x"87"),
   783 => (x"30",x"c1",x"48",x"66"),
   784 => (x"6e",x"58",x"a6",x"d4"),
   785 => (x"70",x"30",x"c1",x"48"),
   786 => (x"48",x"66",x"d4",x"7e"),
   787 => (x"a6",x"d8",x"80",x"c1"),
   788 => (x"b7",x"e0",x"c0",x"58"),
   789 => (x"f7",x"f8",x"04",x"a8"),
   790 => (x"4c",x"66",x"cc",x"87"),
   791 => (x"b7",x"c2",x"84",x"c1"),
   792 => (x"df",x"f7",x"04",x"ac"),
   793 => (x"c6",x"cd",x"c3",x"87"),
   794 => (x"78",x"66",x"c4",x"48"),
   795 => (x"26",x"8e",x"d8",x"ff"),
   796 => (x"26",x"4c",x"26",x"4d"),
   797 => (x"00",x"4f",x"26",x"4b"),
   798 => (x"1e",x"00",x"00",x"00"),
   799 => (x"49",x"72",x"4a",x"c0"),
   800 => (x"cd",x"c3",x"91",x"c4"),
   801 => (x"79",x"ff",x"81",x"d2"),
   802 => (x"b7",x"c6",x"82",x"c1"),
   803 => (x"87",x"ee",x"04",x"aa"),
   804 => (x"48",x"c6",x"cd",x"c3"),
   805 => (x"78",x"40",x"40",x"c0"),
   806 => (x"73",x"1e",x"4f",x"26"),
   807 => (x"f4",x"4b",x"71",x"1e"),
   808 => (x"49",x"73",x"87",x"c4"),
   809 => (x"87",x"ec",x"f9",x"fe"),
   810 => (x"1e",x"87",x"c8",x"ff"),
   811 => (x"4b",x"c0",x"1e",x"73"),
   812 => (x"49",x"c8",x"f3",x"c2"),
   813 => (x"70",x"87",x"ce",x"ed"),
   814 => (x"87",x"c4",x"05",x"98"),
   815 => (x"4b",x"d4",x"f3",x"c2"),
   816 => (x"73",x"87",x"f8",x"fe"),
   817 => (x"87",x"eb",x"fe",x"48"),
   818 => (x"43",x"49",x"52",x"4f"),
   819 => (x"20",x"20",x"20",x"20"),
   820 => (x"00",x"4d",x"4f",x"52"),
   821 => (x"20",x"4d",x"4f",x"52"),
   822 => (x"64",x"61",x"6f",x"6c"),
   823 => (x"20",x"67",x"6e",x"69"),
   824 => (x"6c",x"69",x"61",x"66"),
   825 => (x"f4",x"00",x"64",x"65"),
   826 => (x"05",x"f5",x"f2",x"eb"),
   827 => (x"03",x"0c",x"04",x"06"),
   828 => (x"66",x"0a",x"83",x"0b"),
   829 => (x"5a",x"00",x"fc",x"00"),
   830 => (x"00",x"00",x"da",x"00"),
   831 => (x"05",x"08",x"94",x"80"),
   832 => (x"02",x"00",x"78",x"80"),
   833 => (x"03",x"00",x"01",x"80"),
   834 => (x"04",x"00",x"09",x"80"),
   835 => (x"01",x"00",x"00",x"80"),
   836 => (x"26",x"08",x"91",x"80"),
   837 => (x"1d",x"00",x"04",x"00"),
   838 => (x"1c",x"00",x"00",x"00"),
   839 => (x"25",x"00",x"00",x"00"),
   840 => (x"1a",x"00",x"0c",x"00"),
   841 => (x"1b",x"00",x"00",x"00"),
   842 => (x"24",x"00",x"00",x"00"),
   843 => (x"12",x"00",x"00",x"00"),
   844 => (x"2e",x"00",x"00",x"01"),
   845 => (x"2d",x"00",x"03",x"00"),
   846 => (x"23",x"00",x"00",x"00"),
   847 => (x"36",x"00",x"00",x"00"),
   848 => (x"21",x"00",x"0b",x"00"),
   849 => (x"2b",x"00",x"00",x"00"),
   850 => (x"2c",x"00",x"00",x"00"),
   851 => (x"22",x"00",x"00",x"00"),
   852 => (x"3d",x"00",x"00",x"00"),
   853 => (x"35",x"00",x"6c",x"00"),
   854 => (x"34",x"00",x"00",x"00"),
   855 => (x"3e",x"00",x"00",x"00"),
   856 => (x"32",x"00",x"75",x"00"),
   857 => (x"33",x"00",x"00",x"00"),
   858 => (x"3c",x"00",x"00",x"00"),
   859 => (x"2a",x"00",x"6b",x"00"),
   860 => (x"46",x"00",x"00",x"00"),
   861 => (x"43",x"00",x"01",x"00"),
   862 => (x"3b",x"00",x"73",x"00"),
   863 => (x"45",x"00",x"69",x"00"),
   864 => (x"3a",x"00",x"09",x"00"),
   865 => (x"42",x"00",x"70",x"00"),
   866 => (x"44",x"00",x"72",x"00"),
   867 => (x"31",x"00",x"74",x"00"),
   868 => (x"55",x"00",x"00",x"00"),
   869 => (x"4d",x"00",x"00",x"00"),
   870 => (x"4b",x"00",x"7c",x"00"),
   871 => (x"7b",x"00",x"7a",x"00"),
   872 => (x"49",x"00",x"00",x"00"),
   873 => (x"4c",x"00",x"71",x"00"),
   874 => (x"54",x"00",x"84",x"00"),
   875 => (x"41",x"00",x"77",x"00"),
   876 => (x"61",x"00",x"00",x"00"),
   877 => (x"5b",x"00",x"00",x"00"),
   878 => (x"52",x"00",x"7c",x"00"),
   879 => (x"f1",x"00",x"00",x"00"),
   880 => (x"59",x"00",x"00",x"00"),
   881 => (x"0e",x"00",x"00",x"02"),
   882 => (x"5d",x"00",x"5d",x"00"),
   883 => (x"4a",x"00",x"00",x"00"),
   884 => (x"16",x"00",x"79",x"00"),
   885 => (x"76",x"00",x"05",x"00"),
   886 => (x"0d",x"00",x"07",x"00"),
   887 => (x"1e",x"00",x"0d",x"00"),
   888 => (x"29",x"00",x"06",x"00"),
   889 => (x"14",x"00",x"00",x"00"),
   890 => (x"15",x"00",x"00",x"04"),
   891 => (x"00",x"00",x"00",x"00"),
   892 => (x"00",x"00",x"00",x"40"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

