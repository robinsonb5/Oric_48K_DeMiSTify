
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"ec",x"cd",x"c3",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"ec",x"cd",x"c3"),
    14 => (x"48",x"f4",x"f7",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"c8",x"e3"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"1e",x"73",x"1e",x"4f"),
    50 => (x"c0",x"02",x"9a",x"72"),
    51 => (x"48",x"c0",x"87",x"e7"),
    52 => (x"a9",x"72",x"4b",x"c1"),
    53 => (x"72",x"87",x"d1",x"06"),
    54 => (x"87",x"c9",x"06",x"82"),
    55 => (x"a9",x"72",x"83",x"73"),
    56 => (x"c3",x"87",x"f4",x"01"),
    57 => (x"3a",x"b2",x"c1",x"87"),
    58 => (x"89",x"03",x"a9",x"72"),
    59 => (x"c1",x"07",x"80",x"73"),
    60 => (x"f3",x"05",x"2b",x"2a"),
    61 => (x"26",x"4b",x"26",x"87"),
    62 => (x"1e",x"75",x"1e",x"4f"),
    63 => (x"b7",x"71",x"4d",x"c4"),
    64 => (x"b9",x"ff",x"04",x"a1"),
    65 => (x"bd",x"c3",x"81",x"c1"),
    66 => (x"a2",x"b7",x"72",x"07"),
    67 => (x"c1",x"ba",x"ff",x"04"),
    68 => (x"07",x"bd",x"c1",x"82"),
    69 => (x"c1",x"87",x"ee",x"fe"),
    70 => (x"b8",x"ff",x"04",x"2d"),
    71 => (x"2d",x"07",x"80",x"c1"),
    72 => (x"c1",x"b9",x"ff",x"04"),
    73 => (x"4d",x"26",x"07",x"81"),
    74 => (x"11",x"1e",x"4f",x"26"),
    75 => (x"08",x"d4",x"ff",x"48"),
    76 => (x"48",x"66",x"c4",x"78"),
    77 => (x"a6",x"c8",x"88",x"c1"),
    78 => (x"05",x"98",x"70",x"58"),
    79 => (x"4f",x"26",x"87",x"ed"),
    80 => (x"48",x"d4",x"ff",x"1e"),
    81 => (x"68",x"78",x"ff",x"c3"),
    82 => (x"48",x"66",x"c4",x"51"),
    83 => (x"a6",x"c8",x"88",x"c1"),
    84 => (x"05",x"98",x"70",x"58"),
    85 => (x"4f",x"26",x"87",x"eb"),
    86 => (x"ff",x"1e",x"73",x"1e"),
    87 => (x"ff",x"c3",x"4b",x"d4"),
    88 => (x"c3",x"4a",x"6b",x"7b"),
    89 => (x"49",x"6b",x"7b",x"ff"),
    90 => (x"b1",x"72",x"32",x"c8"),
    91 => (x"6b",x"7b",x"ff",x"c3"),
    92 => (x"71",x"31",x"c8",x"4a"),
    93 => (x"7b",x"ff",x"c3",x"b2"),
    94 => (x"32",x"c8",x"49",x"6b"),
    95 => (x"48",x"71",x"b1",x"72"),
    96 => (x"4d",x"26",x"87",x"c4"),
    97 => (x"4b",x"26",x"4c",x"26"),
    98 => (x"5e",x"0e",x"4f",x"26"),
    99 => (x"0e",x"5d",x"5c",x"5b"),
   100 => (x"d4",x"ff",x"4a",x"71"),
   101 => (x"c3",x"49",x"72",x"4c"),
   102 => (x"7c",x"71",x"99",x"ff"),
   103 => (x"bf",x"f4",x"f7",x"c2"),
   104 => (x"d0",x"87",x"c8",x"05"),
   105 => (x"30",x"c9",x"48",x"66"),
   106 => (x"d0",x"58",x"a6",x"d4"),
   107 => (x"29",x"d8",x"49",x"66"),
   108 => (x"71",x"99",x"ff",x"c3"),
   109 => (x"49",x"66",x"d0",x"7c"),
   110 => (x"ff",x"c3",x"29",x"d0"),
   111 => (x"d0",x"7c",x"71",x"99"),
   112 => (x"29",x"c8",x"49",x"66"),
   113 => (x"71",x"99",x"ff",x"c3"),
   114 => (x"49",x"66",x"d0",x"7c"),
   115 => (x"71",x"99",x"ff",x"c3"),
   116 => (x"d0",x"49",x"72",x"7c"),
   117 => (x"99",x"ff",x"c3",x"29"),
   118 => (x"4b",x"6c",x"7c",x"71"),
   119 => (x"4d",x"ff",x"f0",x"c9"),
   120 => (x"05",x"ab",x"ff",x"c3"),
   121 => (x"ff",x"c3",x"87",x"d0"),
   122 => (x"c1",x"4b",x"6c",x"7c"),
   123 => (x"87",x"c6",x"02",x"8d"),
   124 => (x"02",x"ab",x"ff",x"c3"),
   125 => (x"48",x"73",x"87",x"f0"),
   126 => (x"1e",x"87",x"c7",x"fe"),
   127 => (x"d4",x"ff",x"49",x"c0"),
   128 => (x"78",x"ff",x"c3",x"48"),
   129 => (x"c8",x"c3",x"81",x"c1"),
   130 => (x"f1",x"04",x"a9",x"b7"),
   131 => (x"1e",x"4f",x"26",x"87"),
   132 => (x"87",x"e7",x"1e",x"73"),
   133 => (x"4b",x"df",x"f8",x"c4"),
   134 => (x"ff",x"c0",x"1e",x"c0"),
   135 => (x"49",x"f7",x"c1",x"f0"),
   136 => (x"c4",x"87",x"e7",x"fd"),
   137 => (x"05",x"a8",x"c1",x"86"),
   138 => (x"ff",x"87",x"ea",x"c0"),
   139 => (x"ff",x"c3",x"48",x"d4"),
   140 => (x"c0",x"c0",x"c1",x"78"),
   141 => (x"1e",x"c0",x"c0",x"c0"),
   142 => (x"c1",x"f0",x"e1",x"c0"),
   143 => (x"c9",x"fd",x"49",x"e9"),
   144 => (x"70",x"86",x"c4",x"87"),
   145 => (x"87",x"ca",x"05",x"98"),
   146 => (x"c3",x"48",x"d4",x"ff"),
   147 => (x"48",x"c1",x"78",x"ff"),
   148 => (x"e6",x"fe",x"87",x"cb"),
   149 => (x"05",x"8b",x"c1",x"87"),
   150 => (x"c0",x"87",x"fd",x"fe"),
   151 => (x"87",x"e6",x"fc",x"48"),
   152 => (x"ff",x"1e",x"73",x"1e"),
   153 => (x"ff",x"c3",x"48",x"d4"),
   154 => (x"c0",x"4b",x"d3",x"78"),
   155 => (x"f0",x"ff",x"c0",x"1e"),
   156 => (x"fc",x"49",x"c1",x"c1"),
   157 => (x"86",x"c4",x"87",x"d4"),
   158 => (x"ca",x"05",x"98",x"70"),
   159 => (x"48",x"d4",x"ff",x"87"),
   160 => (x"c1",x"78",x"ff",x"c3"),
   161 => (x"fd",x"87",x"cb",x"48"),
   162 => (x"8b",x"c1",x"87",x"f1"),
   163 => (x"87",x"db",x"ff",x"05"),
   164 => (x"f1",x"fb",x"48",x"c0"),
   165 => (x"5b",x"5e",x"0e",x"87"),
   166 => (x"d4",x"ff",x"0e",x"5c"),
   167 => (x"87",x"db",x"fd",x"4c"),
   168 => (x"c0",x"1e",x"ea",x"c6"),
   169 => (x"c8",x"c1",x"f0",x"e1"),
   170 => (x"87",x"de",x"fb",x"49"),
   171 => (x"a8",x"c1",x"86",x"c4"),
   172 => (x"fe",x"87",x"c8",x"02"),
   173 => (x"48",x"c0",x"87",x"ea"),
   174 => (x"fa",x"87",x"e2",x"c1"),
   175 => (x"49",x"70",x"87",x"da"),
   176 => (x"99",x"ff",x"ff",x"cf"),
   177 => (x"02",x"a9",x"ea",x"c6"),
   178 => (x"d3",x"fe",x"87",x"c8"),
   179 => (x"c1",x"48",x"c0",x"87"),
   180 => (x"ff",x"c3",x"87",x"cb"),
   181 => (x"4b",x"f1",x"c0",x"7c"),
   182 => (x"70",x"87",x"f4",x"fc"),
   183 => (x"eb",x"c0",x"02",x"98"),
   184 => (x"c0",x"1e",x"c0",x"87"),
   185 => (x"fa",x"c1",x"f0",x"ff"),
   186 => (x"87",x"de",x"fa",x"49"),
   187 => (x"98",x"70",x"86",x"c4"),
   188 => (x"c3",x"87",x"d9",x"05"),
   189 => (x"49",x"6c",x"7c",x"ff"),
   190 => (x"7c",x"7c",x"ff",x"c3"),
   191 => (x"c0",x"c1",x"7c",x"7c"),
   192 => (x"87",x"c4",x"02",x"99"),
   193 => (x"87",x"d5",x"48",x"c1"),
   194 => (x"87",x"d1",x"48",x"c0"),
   195 => (x"c4",x"05",x"ab",x"c2"),
   196 => (x"c8",x"48",x"c0",x"87"),
   197 => (x"05",x"8b",x"c1",x"87"),
   198 => (x"c0",x"87",x"fd",x"fe"),
   199 => (x"87",x"e4",x"f9",x"48"),
   200 => (x"c2",x"1e",x"73",x"1e"),
   201 => (x"c1",x"48",x"f4",x"f7"),
   202 => (x"ff",x"4b",x"c7",x"78"),
   203 => (x"78",x"c2",x"48",x"d0"),
   204 => (x"ff",x"87",x"c8",x"fb"),
   205 => (x"78",x"c3",x"48",x"d0"),
   206 => (x"e5",x"c0",x"1e",x"c0"),
   207 => (x"49",x"c0",x"c1",x"d0"),
   208 => (x"c4",x"87",x"c7",x"f9"),
   209 => (x"05",x"a8",x"c1",x"86"),
   210 => (x"c2",x"4b",x"87",x"c1"),
   211 => (x"87",x"c5",x"05",x"ab"),
   212 => (x"f9",x"c0",x"48",x"c0"),
   213 => (x"05",x"8b",x"c1",x"87"),
   214 => (x"fc",x"87",x"d0",x"ff"),
   215 => (x"f7",x"c2",x"87",x"f7"),
   216 => (x"98",x"70",x"58",x"f8"),
   217 => (x"c1",x"87",x"cd",x"05"),
   218 => (x"f0",x"ff",x"c0",x"1e"),
   219 => (x"f8",x"49",x"d0",x"c1"),
   220 => (x"86",x"c4",x"87",x"d8"),
   221 => (x"c3",x"48",x"d4",x"ff"),
   222 => (x"e0",x"c4",x"78",x"ff"),
   223 => (x"fc",x"f7",x"c2",x"87"),
   224 => (x"48",x"d0",x"ff",x"58"),
   225 => (x"d4",x"ff",x"78",x"c2"),
   226 => (x"78",x"ff",x"c3",x"48"),
   227 => (x"f5",x"f7",x"48",x"c1"),
   228 => (x"5b",x"5e",x"0e",x"87"),
   229 => (x"71",x"0e",x"5d",x"5c"),
   230 => (x"4d",x"ff",x"c3",x"4a"),
   231 => (x"75",x"4c",x"d4",x"ff"),
   232 => (x"48",x"d0",x"ff",x"7c"),
   233 => (x"75",x"78",x"c3",x"c4"),
   234 => (x"c0",x"1e",x"72",x"7c"),
   235 => (x"d8",x"c1",x"f0",x"ff"),
   236 => (x"87",x"d6",x"f7",x"49"),
   237 => (x"98",x"70",x"86",x"c4"),
   238 => (x"c0",x"87",x"c5",x"02"),
   239 => (x"87",x"f0",x"c0",x"48"),
   240 => (x"fe",x"c3",x"7c",x"75"),
   241 => (x"1e",x"c0",x"c8",x"7c"),
   242 => (x"f5",x"49",x"66",x"d4"),
   243 => (x"86",x"c4",x"87",x"dc"),
   244 => (x"7c",x"75",x"7c",x"75"),
   245 => (x"da",x"d8",x"7c",x"75"),
   246 => (x"7c",x"75",x"4b",x"e0"),
   247 => (x"05",x"99",x"49",x"6c"),
   248 => (x"8b",x"c1",x"87",x"c5"),
   249 => (x"75",x"87",x"f3",x"05"),
   250 => (x"48",x"d0",x"ff",x"7c"),
   251 => (x"48",x"c1",x"78",x"c2"),
   252 => (x"1e",x"87",x"cf",x"f6"),
   253 => (x"ff",x"4a",x"d4",x"ff"),
   254 => (x"d1",x"c4",x"48",x"d0"),
   255 => (x"7a",x"ff",x"c3",x"78"),
   256 => (x"f8",x"05",x"89",x"c1"),
   257 => (x"1e",x"4f",x"26",x"87"),
   258 => (x"4b",x"71",x"1e",x"73"),
   259 => (x"df",x"cd",x"ee",x"c5"),
   260 => (x"48",x"d4",x"ff",x"4a"),
   261 => (x"68",x"78",x"ff",x"c3"),
   262 => (x"a8",x"fe",x"c3",x"48"),
   263 => (x"c1",x"87",x"c5",x"02"),
   264 => (x"87",x"ed",x"05",x"8a"),
   265 => (x"c5",x"05",x"9a",x"72"),
   266 => (x"c0",x"48",x"c0",x"87"),
   267 => (x"9b",x"73",x"87",x"ea"),
   268 => (x"c8",x"87",x"cc",x"02"),
   269 => (x"49",x"73",x"1e",x"66"),
   270 => (x"c4",x"87",x"c5",x"f4"),
   271 => (x"c8",x"87",x"c6",x"86"),
   272 => (x"ee",x"fe",x"49",x"66"),
   273 => (x"48",x"d4",x"ff",x"87"),
   274 => (x"78",x"78",x"ff",x"c3"),
   275 => (x"c5",x"05",x"9b",x"73"),
   276 => (x"48",x"d0",x"ff",x"87"),
   277 => (x"48",x"c1",x"78",x"d0"),
   278 => (x"1e",x"87",x"eb",x"f4"),
   279 => (x"4a",x"71",x"1e",x"73"),
   280 => (x"d4",x"ff",x"4b",x"c0"),
   281 => (x"78",x"ff",x"c3",x"48"),
   282 => (x"c4",x"48",x"d0",x"ff"),
   283 => (x"d4",x"ff",x"78",x"c3"),
   284 => (x"78",x"ff",x"c3",x"48"),
   285 => (x"ff",x"c0",x"1e",x"72"),
   286 => (x"49",x"d1",x"c1",x"f0"),
   287 => (x"c4",x"87",x"cb",x"f4"),
   288 => (x"05",x"98",x"70",x"86"),
   289 => (x"c0",x"c8",x"87",x"cd"),
   290 => (x"49",x"66",x"cc",x"1e"),
   291 => (x"c4",x"87",x"f8",x"fd"),
   292 => (x"ff",x"4b",x"70",x"86"),
   293 => (x"78",x"c2",x"48",x"d0"),
   294 => (x"e9",x"f3",x"48",x"73"),
   295 => (x"5b",x"5e",x"0e",x"87"),
   296 => (x"c0",x"0e",x"5d",x"5c"),
   297 => (x"f0",x"ff",x"c0",x"1e"),
   298 => (x"f3",x"49",x"c9",x"c1"),
   299 => (x"1e",x"d2",x"87",x"dc"),
   300 => (x"49",x"fc",x"f7",x"c2"),
   301 => (x"c8",x"87",x"d0",x"fd"),
   302 => (x"c1",x"4c",x"c0",x"86"),
   303 => (x"ac",x"b7",x"d2",x"84"),
   304 => (x"c2",x"87",x"f8",x"04"),
   305 => (x"bf",x"97",x"fc",x"f7"),
   306 => (x"99",x"c0",x"c3",x"49"),
   307 => (x"05",x"a9",x"c0",x"c1"),
   308 => (x"c2",x"87",x"e7",x"c0"),
   309 => (x"bf",x"97",x"c3",x"f8"),
   310 => (x"c2",x"31",x"d0",x"49"),
   311 => (x"bf",x"97",x"c4",x"f8"),
   312 => (x"72",x"32",x"c8",x"4a"),
   313 => (x"c5",x"f8",x"c2",x"b1"),
   314 => (x"b1",x"4a",x"bf",x"97"),
   315 => (x"ff",x"cf",x"4c",x"71"),
   316 => (x"c1",x"9c",x"ff",x"ff"),
   317 => (x"c1",x"34",x"ca",x"84"),
   318 => (x"f8",x"c2",x"87",x"e7"),
   319 => (x"49",x"bf",x"97",x"c5"),
   320 => (x"99",x"c6",x"31",x"c1"),
   321 => (x"97",x"c6",x"f8",x"c2"),
   322 => (x"b7",x"c7",x"4a",x"bf"),
   323 => (x"c2",x"b1",x"72",x"2a"),
   324 => (x"bf",x"97",x"c1",x"f8"),
   325 => (x"9d",x"cf",x"4d",x"4a"),
   326 => (x"97",x"c2",x"f8",x"c2"),
   327 => (x"9a",x"c3",x"4a",x"bf"),
   328 => (x"f8",x"c2",x"32",x"ca"),
   329 => (x"4b",x"bf",x"97",x"c3"),
   330 => (x"b2",x"73",x"33",x"c2"),
   331 => (x"97",x"c4",x"f8",x"c2"),
   332 => (x"c0",x"c3",x"4b",x"bf"),
   333 => (x"2b",x"b7",x"c6",x"9b"),
   334 => (x"81",x"c2",x"b2",x"73"),
   335 => (x"30",x"71",x"48",x"c1"),
   336 => (x"48",x"c1",x"49",x"70"),
   337 => (x"4d",x"70",x"30",x"75"),
   338 => (x"84",x"c1",x"4c",x"72"),
   339 => (x"c0",x"c8",x"94",x"71"),
   340 => (x"cc",x"06",x"ad",x"b7"),
   341 => (x"b7",x"34",x"c1",x"87"),
   342 => (x"b7",x"c0",x"c8",x"2d"),
   343 => (x"f4",x"ff",x"01",x"ad"),
   344 => (x"f0",x"48",x"74",x"87"),
   345 => (x"5e",x"0e",x"87",x"dc"),
   346 => (x"0e",x"5d",x"5c",x"5b"),
   347 => (x"c0",x"c3",x"86",x"f8"),
   348 => (x"78",x"c0",x"48",x"e2"),
   349 => (x"1e",x"da",x"f8",x"c2"),
   350 => (x"de",x"fb",x"49",x"c0"),
   351 => (x"70",x"86",x"c4",x"87"),
   352 => (x"87",x"c5",x"05",x"98"),
   353 => (x"ce",x"c9",x"48",x"c0"),
   354 => (x"c1",x"4d",x"c0",x"87"),
   355 => (x"c1",x"fa",x"c0",x"7e"),
   356 => (x"f9",x"c2",x"49",x"bf"),
   357 => (x"c8",x"71",x"4a",x"d0"),
   358 => (x"87",x"ce",x"eb",x"4b"),
   359 => (x"c2",x"05",x"98",x"70"),
   360 => (x"c0",x"7e",x"c0",x"87"),
   361 => (x"49",x"bf",x"fd",x"f9"),
   362 => (x"4a",x"ec",x"f9",x"c2"),
   363 => (x"ea",x"4b",x"c8",x"71"),
   364 => (x"98",x"70",x"87",x"f8"),
   365 => (x"c0",x"87",x"c2",x"05"),
   366 => (x"c0",x"02",x"6e",x"7e"),
   367 => (x"ff",x"c2",x"87",x"fd"),
   368 => (x"c3",x"4d",x"bf",x"e0"),
   369 => (x"bf",x"9f",x"d8",x"c0"),
   370 => (x"d6",x"c5",x"48",x"7e"),
   371 => (x"c7",x"05",x"a8",x"ea"),
   372 => (x"e0",x"ff",x"c2",x"87"),
   373 => (x"87",x"ce",x"4d",x"bf"),
   374 => (x"e9",x"ca",x"48",x"6e"),
   375 => (x"c5",x"02",x"a8",x"d5"),
   376 => (x"c7",x"48",x"c0",x"87"),
   377 => (x"f8",x"c2",x"87",x"f1"),
   378 => (x"49",x"75",x"1e",x"da"),
   379 => (x"c4",x"87",x"ec",x"f9"),
   380 => (x"05",x"98",x"70",x"86"),
   381 => (x"48",x"c0",x"87",x"c5"),
   382 => (x"c0",x"87",x"dc",x"c7"),
   383 => (x"49",x"bf",x"fd",x"f9"),
   384 => (x"4a",x"ec",x"f9",x"c2"),
   385 => (x"e9",x"4b",x"c8",x"71"),
   386 => (x"98",x"70",x"87",x"e0"),
   387 => (x"c3",x"87",x"c8",x"05"),
   388 => (x"c1",x"48",x"e2",x"c0"),
   389 => (x"c0",x"87",x"da",x"78"),
   390 => (x"49",x"bf",x"c1",x"fa"),
   391 => (x"4a",x"d0",x"f9",x"c2"),
   392 => (x"e9",x"4b",x"c8",x"71"),
   393 => (x"98",x"70",x"87",x"c4"),
   394 => (x"87",x"c5",x"c0",x"02"),
   395 => (x"e6",x"c6",x"48",x"c0"),
   396 => (x"d8",x"c0",x"c3",x"87"),
   397 => (x"c1",x"49",x"bf",x"97"),
   398 => (x"c0",x"05",x"a9",x"d5"),
   399 => (x"c0",x"c3",x"87",x"cd"),
   400 => (x"49",x"bf",x"97",x"d9"),
   401 => (x"02",x"a9",x"ea",x"c2"),
   402 => (x"c0",x"87",x"c5",x"c0"),
   403 => (x"87",x"c7",x"c6",x"48"),
   404 => (x"97",x"da",x"f8",x"c2"),
   405 => (x"c3",x"48",x"7e",x"bf"),
   406 => (x"c0",x"02",x"a8",x"e9"),
   407 => (x"48",x"6e",x"87",x"ce"),
   408 => (x"02",x"a8",x"eb",x"c3"),
   409 => (x"c0",x"87",x"c5",x"c0"),
   410 => (x"87",x"eb",x"c5",x"48"),
   411 => (x"97",x"e5",x"f8",x"c2"),
   412 => (x"05",x"99",x"49",x"bf"),
   413 => (x"c2",x"87",x"cc",x"c0"),
   414 => (x"bf",x"97",x"e6",x"f8"),
   415 => (x"02",x"a9",x"c2",x"49"),
   416 => (x"c0",x"87",x"c5",x"c0"),
   417 => (x"87",x"cf",x"c5",x"48"),
   418 => (x"97",x"e7",x"f8",x"c2"),
   419 => (x"c0",x"c3",x"48",x"bf"),
   420 => (x"4c",x"70",x"58",x"de"),
   421 => (x"c3",x"88",x"c1",x"48"),
   422 => (x"c2",x"58",x"e2",x"c0"),
   423 => (x"bf",x"97",x"e8",x"f8"),
   424 => (x"c2",x"81",x"75",x"49"),
   425 => (x"bf",x"97",x"e9",x"f8"),
   426 => (x"72",x"32",x"c8",x"4a"),
   427 => (x"c4",x"c3",x"7e",x"a1"),
   428 => (x"78",x"6e",x"48",x"ef"),
   429 => (x"97",x"ea",x"f8",x"c2"),
   430 => (x"a6",x"c8",x"48",x"bf"),
   431 => (x"e2",x"c0",x"c3",x"58"),
   432 => (x"d4",x"c2",x"02",x"bf"),
   433 => (x"fd",x"f9",x"c0",x"87"),
   434 => (x"f9",x"c2",x"49",x"bf"),
   435 => (x"c8",x"71",x"4a",x"ec"),
   436 => (x"87",x"d6",x"e6",x"4b"),
   437 => (x"c0",x"02",x"98",x"70"),
   438 => (x"48",x"c0",x"87",x"c5"),
   439 => (x"c3",x"87",x"f8",x"c3"),
   440 => (x"4c",x"bf",x"da",x"c0"),
   441 => (x"5c",x"c3",x"c5",x"c3"),
   442 => (x"97",x"ff",x"f8",x"c2"),
   443 => (x"31",x"c8",x"49",x"bf"),
   444 => (x"97",x"fe",x"f8",x"c2"),
   445 => (x"49",x"a1",x"4a",x"bf"),
   446 => (x"97",x"c0",x"f9",x"c2"),
   447 => (x"32",x"d0",x"4a",x"bf"),
   448 => (x"c2",x"49",x"a1",x"72"),
   449 => (x"bf",x"97",x"c1",x"f9"),
   450 => (x"72",x"32",x"d8",x"4a"),
   451 => (x"66",x"c4",x"49",x"a1"),
   452 => (x"ef",x"c4",x"c3",x"91"),
   453 => (x"c4",x"c3",x"81",x"bf"),
   454 => (x"f9",x"c2",x"59",x"f7"),
   455 => (x"4a",x"bf",x"97",x"c7"),
   456 => (x"f9",x"c2",x"32",x"c8"),
   457 => (x"4b",x"bf",x"97",x"c6"),
   458 => (x"f9",x"c2",x"4a",x"a2"),
   459 => (x"4b",x"bf",x"97",x"c8"),
   460 => (x"a2",x"73",x"33",x"d0"),
   461 => (x"c9",x"f9",x"c2",x"4a"),
   462 => (x"cf",x"4b",x"bf",x"97"),
   463 => (x"73",x"33",x"d8",x"9b"),
   464 => (x"c4",x"c3",x"4a",x"a2"),
   465 => (x"c4",x"c3",x"5a",x"fb"),
   466 => (x"c2",x"4a",x"bf",x"f7"),
   467 => (x"c3",x"92",x"74",x"8a"),
   468 => (x"72",x"48",x"fb",x"c4"),
   469 => (x"ca",x"c1",x"78",x"a1"),
   470 => (x"ec",x"f8",x"c2",x"87"),
   471 => (x"c8",x"49",x"bf",x"97"),
   472 => (x"eb",x"f8",x"c2",x"31"),
   473 => (x"a1",x"4a",x"bf",x"97"),
   474 => (x"ea",x"c0",x"c3",x"49"),
   475 => (x"e6",x"c0",x"c3",x"59"),
   476 => (x"31",x"c5",x"49",x"bf"),
   477 => (x"c9",x"81",x"ff",x"c7"),
   478 => (x"c3",x"c5",x"c3",x"29"),
   479 => (x"f1",x"f8",x"c2",x"59"),
   480 => (x"c8",x"4a",x"bf",x"97"),
   481 => (x"f0",x"f8",x"c2",x"32"),
   482 => (x"a2",x"4b",x"bf",x"97"),
   483 => (x"92",x"66",x"c4",x"4a"),
   484 => (x"c4",x"c3",x"82",x"6e"),
   485 => (x"c4",x"c3",x"5a",x"ff"),
   486 => (x"78",x"c0",x"48",x"f7"),
   487 => (x"48",x"f3",x"c4",x"c3"),
   488 => (x"c3",x"78",x"a1",x"72"),
   489 => (x"c3",x"48",x"c3",x"c5"),
   490 => (x"78",x"bf",x"f7",x"c4"),
   491 => (x"48",x"c7",x"c5",x"c3"),
   492 => (x"bf",x"fb",x"c4",x"c3"),
   493 => (x"e2",x"c0",x"c3",x"78"),
   494 => (x"c9",x"c0",x"02",x"bf"),
   495 => (x"c4",x"48",x"74",x"87"),
   496 => (x"c0",x"7e",x"70",x"30"),
   497 => (x"c4",x"c3",x"87",x"c9"),
   498 => (x"c4",x"48",x"bf",x"ff"),
   499 => (x"c3",x"7e",x"70",x"30"),
   500 => (x"6e",x"48",x"e6",x"c0"),
   501 => (x"f8",x"48",x"c1",x"78"),
   502 => (x"26",x"4d",x"26",x"8e"),
   503 => (x"26",x"4b",x"26",x"4c"),
   504 => (x"5b",x"5e",x"0e",x"4f"),
   505 => (x"71",x"0e",x"5d",x"5c"),
   506 => (x"e2",x"c0",x"c3",x"4a"),
   507 => (x"87",x"cb",x"02",x"bf"),
   508 => (x"2b",x"c7",x"4b",x"72"),
   509 => (x"ff",x"c1",x"4c",x"72"),
   510 => (x"72",x"87",x"c9",x"9c"),
   511 => (x"72",x"2b",x"c8",x"4b"),
   512 => (x"9c",x"ff",x"c3",x"4c"),
   513 => (x"bf",x"ef",x"c4",x"c3"),
   514 => (x"f9",x"f9",x"c0",x"83"),
   515 => (x"d9",x"02",x"ab",x"bf"),
   516 => (x"fd",x"f9",x"c0",x"87"),
   517 => (x"da",x"f8",x"c2",x"5b"),
   518 => (x"f0",x"49",x"73",x"1e"),
   519 => (x"86",x"c4",x"87",x"fd"),
   520 => (x"c5",x"05",x"98",x"70"),
   521 => (x"c0",x"48",x"c0",x"87"),
   522 => (x"c0",x"c3",x"87",x"e6"),
   523 => (x"d2",x"02",x"bf",x"e2"),
   524 => (x"c4",x"49",x"74",x"87"),
   525 => (x"da",x"f8",x"c2",x"91"),
   526 => (x"cf",x"4d",x"69",x"81"),
   527 => (x"ff",x"ff",x"ff",x"ff"),
   528 => (x"74",x"87",x"cb",x"9d"),
   529 => (x"c2",x"91",x"c2",x"49"),
   530 => (x"9f",x"81",x"da",x"f8"),
   531 => (x"48",x"75",x"4d",x"69"),
   532 => (x"0e",x"87",x"c6",x"fe"),
   533 => (x"5d",x"5c",x"5b",x"5e"),
   534 => (x"4d",x"71",x"1e",x"0e"),
   535 => (x"49",x"c1",x"1e",x"c0"),
   536 => (x"c4",x"87",x"fe",x"d0"),
   537 => (x"9c",x"4c",x"70",x"86"),
   538 => (x"87",x"c2",x"c1",x"02"),
   539 => (x"4a",x"ea",x"c0",x"c3"),
   540 => (x"df",x"ff",x"49",x"75"),
   541 => (x"98",x"70",x"87",x"d9"),
   542 => (x"87",x"f2",x"c0",x"02"),
   543 => (x"49",x"75",x"4a",x"74"),
   544 => (x"df",x"ff",x"4b",x"cb"),
   545 => (x"98",x"70",x"87",x"fe"),
   546 => (x"87",x"e2",x"c0",x"02"),
   547 => (x"9c",x"74",x"1e",x"c0"),
   548 => (x"c4",x"87",x"c7",x"02"),
   549 => (x"78",x"c0",x"48",x"a6"),
   550 => (x"a6",x"c4",x"87",x"c5"),
   551 => (x"c4",x"78",x"c1",x"48"),
   552 => (x"fc",x"cf",x"49",x"66"),
   553 => (x"70",x"86",x"c4",x"87"),
   554 => (x"fe",x"05",x"9c",x"4c"),
   555 => (x"48",x"74",x"87",x"fe"),
   556 => (x"87",x"e5",x"fc",x"26"),
   557 => (x"5c",x"5b",x"5e",x"0e"),
   558 => (x"86",x"f8",x"0e",x"5d"),
   559 => (x"05",x"9b",x"4b",x"71"),
   560 => (x"48",x"c0",x"87",x"c5"),
   561 => (x"c8",x"87",x"dd",x"c2"),
   562 => (x"7d",x"c0",x"4d",x"a3"),
   563 => (x"c7",x"02",x"66",x"d8"),
   564 => (x"97",x"66",x"d8",x"87"),
   565 => (x"87",x"c5",x"05",x"bf"),
   566 => (x"c7",x"c2",x"48",x"c0"),
   567 => (x"49",x"66",x"d8",x"87"),
   568 => (x"70",x"87",x"f0",x"fd"),
   569 => (x"c1",x"02",x"6e",x"7e"),
   570 => (x"49",x"6e",x"87",x"f8"),
   571 => (x"7d",x"69",x"81",x"dc"),
   572 => (x"81",x"da",x"49",x"6e"),
   573 => (x"9f",x"4c",x"a3",x"c4"),
   574 => (x"c0",x"c3",x"7c",x"69"),
   575 => (x"d0",x"02",x"bf",x"e2"),
   576 => (x"d4",x"49",x"6e",x"87"),
   577 => (x"49",x"69",x"9f",x"81"),
   578 => (x"ff",x"ff",x"c0",x"4a"),
   579 => (x"c2",x"32",x"d0",x"9a"),
   580 => (x"72",x"4a",x"c0",x"87"),
   581 => (x"80",x"6c",x"48",x"49"),
   582 => (x"7b",x"c0",x"7c",x"70"),
   583 => (x"6c",x"49",x"a3",x"cc"),
   584 => (x"49",x"a3",x"d0",x"79"),
   585 => (x"a6",x"c4",x"79",x"c0"),
   586 => (x"d4",x"78",x"c0",x"48"),
   587 => (x"66",x"c4",x"4a",x"a3"),
   588 => (x"72",x"91",x"c8",x"49"),
   589 => (x"41",x"c0",x"49",x"a1"),
   590 => (x"66",x"c4",x"79",x"6c"),
   591 => (x"c8",x"80",x"c1",x"48"),
   592 => (x"b7",x"c6",x"58",x"a6"),
   593 => (x"e2",x"ff",x"04",x"a8"),
   594 => (x"c9",x"4a",x"6d",x"87"),
   595 => (x"c0",x"49",x"72",x"2a"),
   596 => (x"dd",x"ff",x"4a",x"f0"),
   597 => (x"4a",x"70",x"87",x"ef"),
   598 => (x"49",x"a3",x"c4",x"c1"),
   599 => (x"48",x"6e",x"79",x"72"),
   600 => (x"48",x"c0",x"87",x"c2"),
   601 => (x"f0",x"f9",x"8e",x"f8"),
   602 => (x"5b",x"5e",x"0e",x"87"),
   603 => (x"71",x"0e",x"5d",x"5c"),
   604 => (x"f9",x"f9",x"c0",x"4c"),
   605 => (x"74",x"78",x"ff",x"48"),
   606 => (x"ca",x"c1",x"02",x"9c"),
   607 => (x"49",x"a4",x"c8",x"87"),
   608 => (x"c2",x"c1",x"02",x"69"),
   609 => (x"4a",x"66",x"d0",x"87"),
   610 => (x"d4",x"82",x"49",x"6c"),
   611 => (x"66",x"d0",x"5a",x"a6"),
   612 => (x"c0",x"c3",x"b9",x"4d"),
   613 => (x"ff",x"4a",x"bf",x"de"),
   614 => (x"71",x"99",x"72",x"ba"),
   615 => (x"e4",x"c0",x"02",x"99"),
   616 => (x"4b",x"a4",x"c4",x"87"),
   617 => (x"f8",x"f8",x"49",x"6b"),
   618 => (x"c3",x"7b",x"70",x"87"),
   619 => (x"49",x"bf",x"da",x"c0"),
   620 => (x"7c",x"71",x"81",x"6c"),
   621 => (x"c0",x"c3",x"b9",x"75"),
   622 => (x"ff",x"4a",x"bf",x"de"),
   623 => (x"71",x"99",x"72",x"ba"),
   624 => (x"dc",x"ff",x"05",x"99"),
   625 => (x"f8",x"7c",x"75",x"87"),
   626 => (x"73",x"1e",x"87",x"cf"),
   627 => (x"9b",x"4b",x"71",x"1e"),
   628 => (x"c8",x"87",x"c7",x"02"),
   629 => (x"05",x"69",x"49",x"a3"),
   630 => (x"48",x"c0",x"87",x"c5"),
   631 => (x"c3",x"87",x"eb",x"c0"),
   632 => (x"4a",x"bf",x"f3",x"c4"),
   633 => (x"69",x"49",x"a3",x"c4"),
   634 => (x"c3",x"89",x"c2",x"49"),
   635 => (x"91",x"bf",x"da",x"c0"),
   636 => (x"c3",x"4a",x"a2",x"71"),
   637 => (x"49",x"bf",x"de",x"c0"),
   638 => (x"a2",x"71",x"99",x"6b"),
   639 => (x"1e",x"66",x"c8",x"4a"),
   640 => (x"d6",x"e9",x"49",x"72"),
   641 => (x"70",x"86",x"c4",x"87"),
   642 => (x"d0",x"f7",x"48",x"49"),
   643 => (x"1e",x"73",x"1e",x"87"),
   644 => (x"02",x"9b",x"4b",x"71"),
   645 => (x"a3",x"c8",x"87",x"c7"),
   646 => (x"c5",x"05",x"69",x"49"),
   647 => (x"c0",x"48",x"c0",x"87"),
   648 => (x"c4",x"c3",x"87",x"eb"),
   649 => (x"c4",x"4a",x"bf",x"f3"),
   650 => (x"49",x"69",x"49",x"a3"),
   651 => (x"c0",x"c3",x"89",x"c2"),
   652 => (x"71",x"91",x"bf",x"da"),
   653 => (x"c0",x"c3",x"4a",x"a2"),
   654 => (x"6b",x"49",x"bf",x"de"),
   655 => (x"4a",x"a2",x"71",x"99"),
   656 => (x"72",x"1e",x"66",x"c8"),
   657 => (x"87",x"c9",x"e5",x"49"),
   658 => (x"49",x"70",x"86",x"c4"),
   659 => (x"87",x"cd",x"f6",x"48"),
   660 => (x"5c",x"5b",x"5e",x"0e"),
   661 => (x"86",x"f8",x"0e",x"5d"),
   662 => (x"a6",x"c4",x"4b",x"71"),
   663 => (x"c8",x"78",x"ff",x"48"),
   664 => (x"4d",x"69",x"49",x"a3"),
   665 => (x"a3",x"d4",x"4c",x"c0"),
   666 => (x"c8",x"49",x"74",x"4a"),
   667 => (x"49",x"a1",x"72",x"91"),
   668 => (x"66",x"d8",x"49",x"69"),
   669 => (x"70",x"88",x"71",x"48"),
   670 => (x"a9",x"66",x"d8",x"7e"),
   671 => (x"6e",x"87",x"ca",x"01"),
   672 => (x"87",x"c5",x"06",x"ad"),
   673 => (x"6e",x"5c",x"a6",x"c8"),
   674 => (x"c6",x"84",x"c1",x"4d"),
   675 => (x"ff",x"04",x"ac",x"b7"),
   676 => (x"66",x"c4",x"87",x"d4"),
   677 => (x"f4",x"8e",x"f8",x"48"),
   678 => (x"5e",x"0e",x"87",x"ff"),
   679 => (x"0e",x"5d",x"5c",x"5b"),
   680 => (x"a6",x"c8",x"86",x"ec"),
   681 => (x"48",x"a6",x"c8",x"59"),
   682 => (x"ff",x"ff",x"ff",x"c1"),
   683 => (x"c4",x"78",x"ff",x"ff"),
   684 => (x"c0",x"78",x"ff",x"80"),
   685 => (x"c4",x"4c",x"c0",x"4d"),
   686 => (x"83",x"d4",x"4b",x"66"),
   687 => (x"91",x"c8",x"49",x"74"),
   688 => (x"75",x"49",x"a1",x"73"),
   689 => (x"73",x"92",x"c8",x"4a"),
   690 => (x"49",x"69",x"7e",x"a2"),
   691 => (x"d4",x"89",x"bf",x"6e"),
   692 => (x"ad",x"74",x"59",x"a6"),
   693 => (x"d0",x"87",x"c6",x"05"),
   694 => (x"bf",x"6e",x"48",x"a6"),
   695 => (x"48",x"66",x"d0",x"78"),
   696 => (x"04",x"a8",x"b7",x"c0"),
   697 => (x"66",x"d0",x"87",x"cf"),
   698 => (x"a9",x"66",x"c8",x"49"),
   699 => (x"d0",x"87",x"c6",x"03"),
   700 => (x"a6",x"cc",x"5c",x"a6"),
   701 => (x"c6",x"84",x"c1",x"59"),
   702 => (x"fe",x"04",x"ac",x"b7"),
   703 => (x"85",x"c1",x"87",x"f9"),
   704 => (x"04",x"ad",x"b7",x"c6"),
   705 => (x"cc",x"87",x"ee",x"fe"),
   706 => (x"8e",x"ec",x"48",x"66"),
   707 => (x"0e",x"87",x"ca",x"f3"),
   708 => (x"5d",x"5c",x"5b",x"5e"),
   709 => (x"71",x"86",x"f0",x"0e"),
   710 => (x"66",x"e0",x"c0",x"4b"),
   711 => (x"73",x"2c",x"c9",x"4c"),
   712 => (x"e1",x"c3",x"02",x"9b"),
   713 => (x"49",x"a3",x"c8",x"87"),
   714 => (x"d9",x"c3",x"02",x"69"),
   715 => (x"49",x"a3",x"d0",x"87"),
   716 => (x"79",x"66",x"e0",x"c0"),
   717 => (x"02",x"ac",x"7e",x"6b"),
   718 => (x"c3",x"87",x"cb",x"c3"),
   719 => (x"49",x"bf",x"de",x"c0"),
   720 => (x"4a",x"71",x"b9",x"ff"),
   721 => (x"48",x"71",x"9a",x"74"),
   722 => (x"a6",x"cc",x"98",x"6e"),
   723 => (x"4d",x"a3",x"c4",x"58"),
   724 => (x"6d",x"48",x"a6",x"c4"),
   725 => (x"aa",x"66",x"c8",x"78"),
   726 => (x"74",x"87",x"c5",x"05"),
   727 => (x"87",x"d1",x"c2",x"7b"),
   728 => (x"49",x"73",x"1e",x"72"),
   729 => (x"c4",x"87",x"e9",x"fb"),
   730 => (x"48",x"7e",x"70",x"86"),
   731 => (x"04",x"a8",x"b7",x"c0"),
   732 => (x"a3",x"d4",x"87",x"d0"),
   733 => (x"c8",x"49",x"6e",x"4a"),
   734 => (x"49",x"a1",x"72",x"91"),
   735 => (x"7d",x"69",x"7b",x"21"),
   736 => (x"7b",x"c0",x"87",x"c7"),
   737 => (x"69",x"49",x"a3",x"cc"),
   738 => (x"1e",x"66",x"c8",x"7d"),
   739 => (x"ff",x"fa",x"49",x"73"),
   740 => (x"70",x"86",x"c4",x"87"),
   741 => (x"a3",x"c4",x"c1",x"7e"),
   742 => (x"48",x"a6",x"cc",x"49"),
   743 => (x"66",x"c8",x"78",x"69"),
   744 => (x"a8",x"66",x"cc",x"48"),
   745 => (x"6e",x"87",x"c9",x"06"),
   746 => (x"a8",x"b7",x"c0",x"48"),
   747 => (x"87",x"e0",x"c0",x"04"),
   748 => (x"b7",x"c0",x"48",x"6e"),
   749 => (x"ec",x"c0",x"04",x"a8"),
   750 => (x"4a",x"a3",x"d4",x"87"),
   751 => (x"91",x"c8",x"49",x"6e"),
   752 => (x"c8",x"49",x"a1",x"72"),
   753 => (x"88",x"69",x"48",x"66"),
   754 => (x"66",x"cc",x"49",x"70"),
   755 => (x"87",x"d5",x"06",x"a9"),
   756 => (x"c5",x"fb",x"49",x"73"),
   757 => (x"d4",x"49",x"70",x"87"),
   758 => (x"91",x"c8",x"4a",x"a3"),
   759 => (x"c8",x"49",x"a1",x"72"),
   760 => (x"66",x"c4",x"41",x"66"),
   761 => (x"74",x"8c",x"6b",x"79"),
   762 => (x"49",x"73",x"1e",x"49"),
   763 => (x"c4",x"87",x"fa",x"f5"),
   764 => (x"66",x"e0",x"c0",x"86"),
   765 => (x"99",x"ff",x"c7",x"49"),
   766 => (x"c2",x"87",x"cb",x"02"),
   767 => (x"73",x"1e",x"da",x"f8"),
   768 => (x"87",x"c6",x"f7",x"49"),
   769 => (x"8e",x"f0",x"86",x"c4"),
   770 => (x"1e",x"87",x"ce",x"ef"),
   771 => (x"4b",x"71",x"1e",x"73"),
   772 => (x"e4",x"c0",x"02",x"9b"),
   773 => (x"c7",x"c5",x"c3",x"87"),
   774 => (x"c2",x"4a",x"73",x"5b"),
   775 => (x"da",x"c0",x"c3",x"8a"),
   776 => (x"c3",x"92",x"49",x"bf"),
   777 => (x"48",x"bf",x"f3",x"c4"),
   778 => (x"c5",x"c3",x"80",x"72"),
   779 => (x"48",x"71",x"58",x"cb"),
   780 => (x"c0",x"c3",x"30",x"c4"),
   781 => (x"ed",x"c0",x"58",x"ea"),
   782 => (x"c3",x"c5",x"c3",x"87"),
   783 => (x"f7",x"c4",x"c3",x"48"),
   784 => (x"c5",x"c3",x"78",x"bf"),
   785 => (x"c4",x"c3",x"48",x"c7"),
   786 => (x"c3",x"78",x"bf",x"fb"),
   787 => (x"02",x"bf",x"e2",x"c0"),
   788 => (x"c0",x"c3",x"87",x"c9"),
   789 => (x"c4",x"49",x"bf",x"da"),
   790 => (x"c3",x"87",x"c7",x"31"),
   791 => (x"49",x"bf",x"ff",x"c4"),
   792 => (x"c0",x"c3",x"31",x"c4"),
   793 => (x"f4",x"ed",x"59",x"ea"),
   794 => (x"5b",x"5e",x"0e",x"87"),
   795 => (x"4a",x"71",x"0e",x"5c"),
   796 => (x"9a",x"72",x"4b",x"c0"),
   797 => (x"87",x"e1",x"c0",x"02"),
   798 => (x"9f",x"49",x"a2",x"da"),
   799 => (x"c0",x"c3",x"4b",x"69"),
   800 => (x"cf",x"02",x"bf",x"e2"),
   801 => (x"49",x"a2",x"d4",x"87"),
   802 => (x"4c",x"49",x"69",x"9f"),
   803 => (x"9c",x"ff",x"ff",x"c0"),
   804 => (x"87",x"c2",x"34",x"d0"),
   805 => (x"49",x"74",x"4c",x"c0"),
   806 => (x"fd",x"49",x"73",x"b3"),
   807 => (x"fa",x"ec",x"87",x"ed"),
   808 => (x"5b",x"5e",x"0e",x"87"),
   809 => (x"f4",x"0e",x"5d",x"5c"),
   810 => (x"c0",x"4a",x"71",x"86"),
   811 => (x"02",x"9a",x"72",x"7e"),
   812 => (x"f8",x"c2",x"87",x"d8"),
   813 => (x"78",x"c0",x"48",x"d6"),
   814 => (x"48",x"ce",x"f8",x"c2"),
   815 => (x"bf",x"c7",x"c5",x"c3"),
   816 => (x"d2",x"f8",x"c2",x"78"),
   817 => (x"c3",x"c5",x"c3",x"48"),
   818 => (x"c0",x"c3",x"78",x"bf"),
   819 => (x"50",x"c0",x"48",x"f7"),
   820 => (x"bf",x"e6",x"c0",x"c3"),
   821 => (x"d6",x"f8",x"c2",x"49"),
   822 => (x"aa",x"71",x"4a",x"bf"),
   823 => (x"87",x"c0",x"c4",x"03"),
   824 => (x"99",x"cf",x"49",x"72"),
   825 => (x"87",x"e1",x"c0",x"05"),
   826 => (x"1e",x"da",x"f8",x"c2"),
   827 => (x"bf",x"ce",x"f8",x"c2"),
   828 => (x"ce",x"f8",x"c2",x"49"),
   829 => (x"78",x"a1",x"c1",x"48"),
   830 => (x"de",x"dd",x"ff",x"71"),
   831 => (x"c0",x"86",x"c4",x"87"),
   832 => (x"c2",x"48",x"f5",x"f9"),
   833 => (x"cc",x"78",x"da",x"f8"),
   834 => (x"f5",x"f9",x"c0",x"87"),
   835 => (x"e0",x"c0",x"48",x"bf"),
   836 => (x"f9",x"f9",x"c0",x"80"),
   837 => (x"d6",x"f8",x"c2",x"58"),
   838 => (x"80",x"c1",x"48",x"bf"),
   839 => (x"58",x"da",x"f8",x"c2"),
   840 => (x"00",x"0e",x"75",x"27"),
   841 => (x"bf",x"97",x"bf",x"00"),
   842 => (x"c2",x"02",x"9d",x"4d"),
   843 => (x"e5",x"c3",x"87",x"e2"),
   844 => (x"db",x"c2",x"02",x"ad"),
   845 => (x"f5",x"f9",x"c0",x"87"),
   846 => (x"a3",x"cb",x"4b",x"bf"),
   847 => (x"cf",x"4c",x"11",x"49"),
   848 => (x"d2",x"c1",x"05",x"ac"),
   849 => (x"df",x"49",x"75",x"87"),
   850 => (x"cd",x"89",x"c1",x"99"),
   851 => (x"ea",x"c0",x"c3",x"91"),
   852 => (x"4a",x"a3",x"c1",x"81"),
   853 => (x"a3",x"c3",x"51",x"12"),
   854 => (x"c5",x"51",x"12",x"4a"),
   855 => (x"51",x"12",x"4a",x"a3"),
   856 => (x"12",x"4a",x"a3",x"c7"),
   857 => (x"4a",x"a3",x"c9",x"51"),
   858 => (x"a3",x"ce",x"51",x"12"),
   859 => (x"d0",x"51",x"12",x"4a"),
   860 => (x"51",x"12",x"4a",x"a3"),
   861 => (x"12",x"4a",x"a3",x"d2"),
   862 => (x"4a",x"a3",x"d4",x"51"),
   863 => (x"a3",x"d6",x"51",x"12"),
   864 => (x"d8",x"51",x"12",x"4a"),
   865 => (x"51",x"12",x"4a",x"a3"),
   866 => (x"12",x"4a",x"a3",x"dc"),
   867 => (x"4a",x"a3",x"de",x"51"),
   868 => (x"7e",x"c1",x"51",x"12"),
   869 => (x"74",x"87",x"f9",x"c0"),
   870 => (x"05",x"99",x"c8",x"49"),
   871 => (x"74",x"87",x"ea",x"c0"),
   872 => (x"05",x"99",x"d0",x"49"),
   873 => (x"66",x"dc",x"87",x"d0"),
   874 => (x"87",x"ca",x"c0",x"02"),
   875 => (x"66",x"dc",x"49",x"73"),
   876 => (x"02",x"98",x"70",x"0f"),
   877 => (x"05",x"6e",x"87",x"d3"),
   878 => (x"c3",x"87",x"c6",x"c0"),
   879 => (x"c0",x"48",x"ea",x"c0"),
   880 => (x"f5",x"f9",x"c0",x"50"),
   881 => (x"e7",x"c2",x"48",x"bf"),
   882 => (x"f7",x"c0",x"c3",x"87"),
   883 => (x"7e",x"50",x"c0",x"48"),
   884 => (x"bf",x"e6",x"c0",x"c3"),
   885 => (x"d6",x"f8",x"c2",x"49"),
   886 => (x"aa",x"71",x"4a",x"bf"),
   887 => (x"87",x"c0",x"fc",x"04"),
   888 => (x"bf",x"c7",x"c5",x"c3"),
   889 => (x"87",x"c8",x"c0",x"05"),
   890 => (x"bf",x"e2",x"c0",x"c3"),
   891 => (x"87",x"fe",x"c1",x"02"),
   892 => (x"48",x"f9",x"f9",x"c0"),
   893 => (x"f8",x"c2",x"78",x"ff"),
   894 => (x"e7",x"49",x"bf",x"d2"),
   895 => (x"49",x"70",x"87",x"e3"),
   896 => (x"59",x"d6",x"f8",x"c2"),
   897 => (x"c2",x"48",x"a6",x"c4"),
   898 => (x"78",x"bf",x"d2",x"f8"),
   899 => (x"bf",x"e2",x"c0",x"c3"),
   900 => (x"87",x"d8",x"c0",x"02"),
   901 => (x"cf",x"49",x"66",x"c4"),
   902 => (x"f8",x"ff",x"ff",x"ff"),
   903 => (x"c0",x"02",x"a9",x"99"),
   904 => (x"4d",x"c0",x"87",x"c5"),
   905 => (x"c1",x"87",x"e1",x"c0"),
   906 => (x"87",x"dc",x"c0",x"4d"),
   907 => (x"cf",x"49",x"66",x"c4"),
   908 => (x"a9",x"99",x"f8",x"ff"),
   909 => (x"87",x"c8",x"c0",x"02"),
   910 => (x"c0",x"48",x"a6",x"c8"),
   911 => (x"87",x"c5",x"c0",x"78"),
   912 => (x"c1",x"48",x"a6",x"c8"),
   913 => (x"4d",x"66",x"c8",x"78"),
   914 => (x"c0",x"05",x"9d",x"75"),
   915 => (x"66",x"c4",x"87",x"e0"),
   916 => (x"c3",x"89",x"c2",x"49"),
   917 => (x"4a",x"bf",x"da",x"c0"),
   918 => (x"f3",x"c4",x"c3",x"91"),
   919 => (x"f8",x"c2",x"4a",x"bf"),
   920 => (x"a1",x"72",x"48",x"ce"),
   921 => (x"d6",x"f8",x"c2",x"78"),
   922 => (x"f9",x"78",x"c0",x"48"),
   923 => (x"48",x"c0",x"87",x"e2"),
   924 => (x"e4",x"e5",x"8e",x"f4"),
   925 => (x"00",x"00",x"00",x"87"),
   926 => (x"ff",x"ff",x"ff",x"00"),
   927 => (x"00",x"0e",x"85",x"ff"),
   928 => (x"00",x"0e",x"8e",x"00"),
   929 => (x"54",x"41",x"46",x"00"),
   930 => (x"20",x"20",x"32",x"33"),
   931 => (x"41",x"46",x"00",x"20"),
   932 => (x"20",x"36",x"31",x"54"),
   933 => (x"1e",x"00",x"20",x"20"),
   934 => (x"c3",x"48",x"d4",x"ff"),
   935 => (x"48",x"68",x"78",x"ff"),
   936 => (x"ff",x"1e",x"4f",x"26"),
   937 => (x"ff",x"c3",x"48",x"d4"),
   938 => (x"48",x"d0",x"ff",x"78"),
   939 => (x"ff",x"78",x"e1",x"c8"),
   940 => (x"78",x"d4",x"48",x"d4"),
   941 => (x"48",x"cb",x"c5",x"c3"),
   942 => (x"50",x"bf",x"d4",x"ff"),
   943 => (x"ff",x"1e",x"4f",x"26"),
   944 => (x"e0",x"c0",x"48",x"d0"),
   945 => (x"1e",x"4f",x"26",x"78"),
   946 => (x"70",x"87",x"cc",x"ff"),
   947 => (x"c6",x"02",x"99",x"49"),
   948 => (x"a9",x"fb",x"c0",x"87"),
   949 => (x"71",x"87",x"f1",x"05"),
   950 => (x"0e",x"4f",x"26",x"48"),
   951 => (x"0e",x"5c",x"5b",x"5e"),
   952 => (x"4c",x"c0",x"4b",x"71"),
   953 => (x"70",x"87",x"f0",x"fe"),
   954 => (x"c0",x"02",x"99",x"49"),
   955 => (x"ec",x"c0",x"87",x"f9"),
   956 => (x"f2",x"c0",x"02",x"a9"),
   957 => (x"a9",x"fb",x"c0",x"87"),
   958 => (x"87",x"eb",x"c0",x"02"),
   959 => (x"ac",x"b7",x"66",x"cc"),
   960 => (x"d0",x"87",x"c7",x"03"),
   961 => (x"87",x"c2",x"02",x"66"),
   962 => (x"99",x"71",x"53",x"71"),
   963 => (x"c1",x"87",x"c2",x"02"),
   964 => (x"87",x"c3",x"fe",x"84"),
   965 => (x"02",x"99",x"49",x"70"),
   966 => (x"ec",x"c0",x"87",x"cd"),
   967 => (x"87",x"c7",x"02",x"a9"),
   968 => (x"05",x"a9",x"fb",x"c0"),
   969 => (x"d0",x"87",x"d5",x"ff"),
   970 => (x"87",x"c3",x"02",x"66"),
   971 => (x"c0",x"7b",x"97",x"c0"),
   972 => (x"c4",x"05",x"a9",x"ec"),
   973 => (x"c5",x"4a",x"74",x"87"),
   974 => (x"c0",x"4a",x"74",x"87"),
   975 => (x"48",x"72",x"8a",x"0a"),
   976 => (x"4d",x"26",x"87",x"c2"),
   977 => (x"4b",x"26",x"4c",x"26"),
   978 => (x"fd",x"1e",x"4f",x"26"),
   979 => (x"49",x"70",x"87",x"c9"),
   980 => (x"a9",x"b7",x"f0",x"c0"),
   981 => (x"c0",x"87",x"ca",x"04"),
   982 => (x"01",x"a9",x"b7",x"f9"),
   983 => (x"f0",x"c0",x"87",x"c3"),
   984 => (x"b7",x"c1",x"c1",x"89"),
   985 => (x"87",x"ca",x"04",x"a9"),
   986 => (x"a9",x"b7",x"da",x"c1"),
   987 => (x"c0",x"87",x"c3",x"01"),
   988 => (x"48",x"71",x"89",x"f7"),
   989 => (x"5e",x"0e",x"4f",x"26"),
   990 => (x"71",x"0e",x"5c",x"5b"),
   991 => (x"4c",x"d4",x"ff",x"4a"),
   992 => (x"ea",x"c0",x"49",x"72"),
   993 => (x"9b",x"4b",x"70",x"87"),
   994 => (x"c1",x"87",x"c2",x"02"),
   995 => (x"48",x"d0",x"ff",x"8b"),
   996 => (x"c1",x"78",x"c5",x"c8"),
   997 => (x"49",x"73",x"7c",x"d5"),
   998 => (x"e4",x"c2",x"31",x"c6"),
   999 => (x"4a",x"bf",x"97",x"f0"),
  1000 => (x"70",x"b0",x"71",x"48"),
  1001 => (x"48",x"d0",x"ff",x"7c"),
  1002 => (x"48",x"73",x"78",x"c4"),
  1003 => (x"0e",x"87",x"d5",x"fe"),
  1004 => (x"5d",x"5c",x"5b",x"5e"),
  1005 => (x"71",x"86",x"f8",x"0e"),
  1006 => (x"fb",x"7e",x"c0",x"4c"),
  1007 => (x"4b",x"c0",x"87",x"e4"),
  1008 => (x"97",x"dc",x"c1",x"c1"),
  1009 => (x"a9",x"c0",x"49",x"bf"),
  1010 => (x"fb",x"87",x"cf",x"04"),
  1011 => (x"83",x"c1",x"87",x"f9"),
  1012 => (x"97",x"dc",x"c1",x"c1"),
  1013 => (x"06",x"ab",x"49",x"bf"),
  1014 => (x"c1",x"c1",x"87",x"f1"),
  1015 => (x"02",x"bf",x"97",x"dc"),
  1016 => (x"f2",x"fa",x"87",x"cf"),
  1017 => (x"99",x"49",x"70",x"87"),
  1018 => (x"c0",x"87",x"c6",x"02"),
  1019 => (x"f1",x"05",x"a9",x"ec"),
  1020 => (x"fa",x"4b",x"c0",x"87"),
  1021 => (x"4d",x"70",x"87",x"e1"),
  1022 => (x"c8",x"87",x"dc",x"fa"),
  1023 => (x"d6",x"fa",x"58",x"a6"),
  1024 => (x"c1",x"4a",x"70",x"87"),
  1025 => (x"49",x"a4",x"c8",x"83"),
  1026 => (x"ad",x"49",x"69",x"97"),
  1027 => (x"c0",x"87",x"c7",x"02"),
  1028 => (x"c0",x"05",x"ad",x"ff"),
  1029 => (x"a4",x"c9",x"87",x"e7"),
  1030 => (x"49",x"69",x"97",x"49"),
  1031 => (x"02",x"a9",x"66",x"c4"),
  1032 => (x"c0",x"48",x"87",x"c7"),
  1033 => (x"d4",x"05",x"a8",x"ff"),
  1034 => (x"49",x"a4",x"ca",x"87"),
  1035 => (x"aa",x"49",x"69",x"97"),
  1036 => (x"c0",x"87",x"c6",x"02"),
  1037 => (x"c4",x"05",x"aa",x"ff"),
  1038 => (x"d0",x"7e",x"c1",x"87"),
  1039 => (x"ad",x"ec",x"c0",x"87"),
  1040 => (x"c0",x"87",x"c6",x"02"),
  1041 => (x"c4",x"05",x"ad",x"fb"),
  1042 => (x"c1",x"4b",x"c0",x"87"),
  1043 => (x"fe",x"02",x"6e",x"7e"),
  1044 => (x"e9",x"f9",x"87",x"e1"),
  1045 => (x"f8",x"48",x"73",x"87"),
  1046 => (x"87",x"e6",x"fb",x"8e"),
  1047 => (x"5b",x"5e",x"0e",x"00"),
  1048 => (x"1e",x"0e",x"5d",x"5c"),
  1049 => (x"4c",x"c0",x"4b",x"71"),
  1050 => (x"c0",x"04",x"ab",x"4d"),
  1051 => (x"fe",x"c0",x"87",x"e8"),
  1052 => (x"9d",x"75",x"1e",x"ef"),
  1053 => (x"c0",x"87",x"c4",x"02"),
  1054 => (x"c1",x"87",x"c2",x"4a"),
  1055 => (x"f0",x"49",x"72",x"4a"),
  1056 => (x"86",x"c4",x"87",x"df"),
  1057 => (x"84",x"c1",x"7e",x"70"),
  1058 => (x"87",x"c2",x"05",x"6e"),
  1059 => (x"85",x"c1",x"4c",x"73"),
  1060 => (x"ff",x"06",x"ac",x"73"),
  1061 => (x"48",x"6e",x"87",x"d8"),
  1062 => (x"26",x"4d",x"26",x"26"),
  1063 => (x"26",x"4b",x"26",x"4c"),
  1064 => (x"5b",x"5e",x"0e",x"4f"),
  1065 => (x"1e",x"0e",x"5d",x"5c"),
  1066 => (x"de",x"49",x"4c",x"71"),
  1067 => (x"e5",x"c5",x"c3",x"91"),
  1068 => (x"97",x"85",x"71",x"4d"),
  1069 => (x"dd",x"c1",x"02",x"6d"),
  1070 => (x"d0",x"c5",x"c3",x"87"),
  1071 => (x"82",x"74",x"4a",x"bf"),
  1072 => (x"d8",x"fe",x"49",x"72"),
  1073 => (x"6e",x"7e",x"70",x"87"),
  1074 => (x"87",x"f3",x"c0",x"02"),
  1075 => (x"4b",x"d8",x"c5",x"c3"),
  1076 => (x"49",x"cb",x"4a",x"6e"),
  1077 => (x"87",x"d0",x"ff",x"fe"),
  1078 => (x"93",x"cb",x"4b",x"74"),
  1079 => (x"83",x"f7",x"e4",x"c1"),
  1080 => (x"c4",x"c1",x"83",x"c4"),
  1081 => (x"49",x"74",x"7b",x"da"),
  1082 => (x"87",x"d9",x"c2",x"c1"),
  1083 => (x"c5",x"c3",x"7b",x"75"),
  1084 => (x"49",x"bf",x"97",x"e4"),
  1085 => (x"d8",x"c5",x"c3",x"1e"),
  1086 => (x"f5",x"df",x"c1",x"49"),
  1087 => (x"74",x"86",x"c4",x"87"),
  1088 => (x"c0",x"c2",x"c1",x"49"),
  1089 => (x"c1",x"49",x"c0",x"87"),
  1090 => (x"c3",x"87",x"df",x"c3"),
  1091 => (x"c0",x"48",x"cc",x"c5"),
  1092 => (x"dd",x"49",x"c1",x"78"),
  1093 => (x"fd",x"26",x"87",x"cb"),
  1094 => (x"6f",x"4c",x"87",x"ff"),
  1095 => (x"6e",x"69",x"64",x"61"),
  1096 => (x"2e",x"2e",x"2e",x"67"),
  1097 => (x"5b",x"5e",x"0e",x"00"),
  1098 => (x"4b",x"71",x"0e",x"5c"),
  1099 => (x"d0",x"c5",x"c3",x"4a"),
  1100 => (x"49",x"72",x"82",x"bf"),
  1101 => (x"70",x"87",x"e6",x"fc"),
  1102 => (x"c4",x"02",x"9c",x"4c"),
  1103 => (x"e8",x"ec",x"49",x"87"),
  1104 => (x"d0",x"c5",x"c3",x"87"),
  1105 => (x"c1",x"78",x"c0",x"48"),
  1106 => (x"87",x"d5",x"dc",x"49"),
  1107 => (x"0e",x"87",x"cc",x"fd"),
  1108 => (x"5d",x"5c",x"5b",x"5e"),
  1109 => (x"c2",x"86",x"f4",x"0e"),
  1110 => (x"c0",x"4d",x"da",x"f8"),
  1111 => (x"48",x"a6",x"c4",x"4c"),
  1112 => (x"c5",x"c3",x"78",x"c0"),
  1113 => (x"c0",x"49",x"bf",x"d0"),
  1114 => (x"c1",x"c1",x"06",x"a9"),
  1115 => (x"da",x"f8",x"c2",x"87"),
  1116 => (x"c0",x"02",x"98",x"48"),
  1117 => (x"fe",x"c0",x"87",x"f8"),
  1118 => (x"66",x"c8",x"1e",x"ef"),
  1119 => (x"c4",x"87",x"c7",x"02"),
  1120 => (x"78",x"c0",x"48",x"a6"),
  1121 => (x"a6",x"c4",x"87",x"c5"),
  1122 => (x"c4",x"78",x"c1",x"48"),
  1123 => (x"d0",x"ec",x"49",x"66"),
  1124 => (x"70",x"86",x"c4",x"87"),
  1125 => (x"c4",x"84",x"c1",x"4d"),
  1126 => (x"80",x"c1",x"48",x"66"),
  1127 => (x"c3",x"58",x"a6",x"c8"),
  1128 => (x"49",x"bf",x"d0",x"c5"),
  1129 => (x"87",x"c6",x"03",x"ac"),
  1130 => (x"ff",x"05",x"9d",x"75"),
  1131 => (x"4c",x"c0",x"87",x"c8"),
  1132 => (x"c3",x"02",x"9d",x"75"),
  1133 => (x"fe",x"c0",x"87",x"e0"),
  1134 => (x"66",x"c8",x"1e",x"ef"),
  1135 => (x"cc",x"87",x"c7",x"02"),
  1136 => (x"78",x"c0",x"48",x"a6"),
  1137 => (x"a6",x"cc",x"87",x"c5"),
  1138 => (x"cc",x"78",x"c1",x"48"),
  1139 => (x"d0",x"eb",x"49",x"66"),
  1140 => (x"70",x"86",x"c4",x"87"),
  1141 => (x"c2",x"02",x"6e",x"7e"),
  1142 => (x"49",x"6e",x"87",x"e9"),
  1143 => (x"69",x"97",x"81",x"cb"),
  1144 => (x"02",x"99",x"d0",x"49"),
  1145 => (x"c1",x"87",x"d6",x"c1"),
  1146 => (x"74",x"4a",x"e5",x"c4"),
  1147 => (x"c1",x"91",x"cb",x"49"),
  1148 => (x"72",x"81",x"f7",x"e4"),
  1149 => (x"c3",x"81",x"c8",x"79"),
  1150 => (x"49",x"74",x"51",x"ff"),
  1151 => (x"c5",x"c3",x"91",x"de"),
  1152 => (x"85",x"71",x"4d",x"e5"),
  1153 => (x"7d",x"97",x"c1",x"c2"),
  1154 => (x"c0",x"49",x"a5",x"c1"),
  1155 => (x"c0",x"c3",x"51",x"e0"),
  1156 => (x"02",x"bf",x"97",x"ea"),
  1157 => (x"84",x"c1",x"87",x"d2"),
  1158 => (x"c3",x"4b",x"a5",x"c2"),
  1159 => (x"db",x"4a",x"ea",x"c0"),
  1160 => (x"c3",x"fa",x"fe",x"49"),
  1161 => (x"87",x"db",x"c1",x"87"),
  1162 => (x"c0",x"49",x"a5",x"cd"),
  1163 => (x"c2",x"84",x"c1",x"51"),
  1164 => (x"4a",x"6e",x"4b",x"a5"),
  1165 => (x"f9",x"fe",x"49",x"cb"),
  1166 => (x"c6",x"c1",x"87",x"ee"),
  1167 => (x"e1",x"c2",x"c1",x"87"),
  1168 => (x"cb",x"49",x"74",x"4a"),
  1169 => (x"f7",x"e4",x"c1",x"91"),
  1170 => (x"c3",x"79",x"72",x"81"),
  1171 => (x"bf",x"97",x"ea",x"c0"),
  1172 => (x"74",x"87",x"d8",x"02"),
  1173 => (x"c1",x"91",x"de",x"49"),
  1174 => (x"e5",x"c5",x"c3",x"84"),
  1175 => (x"c3",x"83",x"71",x"4b"),
  1176 => (x"dd",x"4a",x"ea",x"c0"),
  1177 => (x"ff",x"f8",x"fe",x"49"),
  1178 => (x"74",x"87",x"d8",x"87"),
  1179 => (x"c3",x"93",x"de",x"4b"),
  1180 => (x"cb",x"83",x"e5",x"c5"),
  1181 => (x"51",x"c0",x"49",x"a3"),
  1182 => (x"6e",x"73",x"84",x"c1"),
  1183 => (x"fe",x"49",x"cb",x"4a"),
  1184 => (x"c4",x"87",x"e5",x"f8"),
  1185 => (x"80",x"c1",x"48",x"66"),
  1186 => (x"c7",x"58",x"a6",x"c8"),
  1187 => (x"c5",x"c0",x"03",x"ac"),
  1188 => (x"fc",x"05",x"6e",x"87"),
  1189 => (x"48",x"74",x"87",x"e0"),
  1190 => (x"fc",x"f7",x"8e",x"f4"),
  1191 => (x"1e",x"73",x"1e",x"87"),
  1192 => (x"cb",x"49",x"4b",x"71"),
  1193 => (x"f7",x"e4",x"c1",x"91"),
  1194 => (x"4a",x"a1",x"c8",x"81"),
  1195 => (x"48",x"f0",x"e4",x"c2"),
  1196 => (x"a1",x"c9",x"50",x"12"),
  1197 => (x"dc",x"c1",x"c1",x"4a"),
  1198 => (x"ca",x"50",x"12",x"48"),
  1199 => (x"e4",x"c5",x"c3",x"81"),
  1200 => (x"c3",x"50",x"11",x"48"),
  1201 => (x"bf",x"97",x"e4",x"c5"),
  1202 => (x"49",x"c0",x"1e",x"49"),
  1203 => (x"87",x"e2",x"d8",x"c1"),
  1204 => (x"48",x"cc",x"c5",x"c3"),
  1205 => (x"49",x"c1",x"78",x"de"),
  1206 => (x"26",x"87",x"c6",x"d6"),
  1207 => (x"1e",x"87",x"fe",x"f6"),
  1208 => (x"cb",x"49",x"4a",x"71"),
  1209 => (x"f7",x"e4",x"c1",x"91"),
  1210 => (x"11",x"81",x"c8",x"81"),
  1211 => (x"d0",x"c5",x"c3",x"48"),
  1212 => (x"d0",x"c5",x"c3",x"58"),
  1213 => (x"c1",x"78",x"c0",x"48"),
  1214 => (x"87",x"e5",x"d5",x"49"),
  1215 => (x"c0",x"1e",x"4f",x"26"),
  1216 => (x"e5",x"fb",x"c0",x"49"),
  1217 => (x"1e",x"4f",x"26",x"87"),
  1218 => (x"d2",x"02",x"99",x"71"),
  1219 => (x"cc",x"e6",x"c1",x"87"),
  1220 => (x"f7",x"50",x"c0",x"48"),
  1221 => (x"df",x"cb",x"c1",x"80"),
  1222 => (x"f0",x"e4",x"c1",x"40"),
  1223 => (x"c1",x"87",x"ce",x"78"),
  1224 => (x"c1",x"48",x"c8",x"e6"),
  1225 => (x"fc",x"78",x"e9",x"e4"),
  1226 => (x"fe",x"cb",x"c1",x"80"),
  1227 => (x"0e",x"4f",x"26",x"78"),
  1228 => (x"0e",x"5c",x"5b",x"5e"),
  1229 => (x"cb",x"4a",x"4c",x"71"),
  1230 => (x"f7",x"e4",x"c1",x"92"),
  1231 => (x"49",x"a2",x"c8",x"82"),
  1232 => (x"97",x"4b",x"a2",x"c9"),
  1233 => (x"97",x"1e",x"4b",x"6b"),
  1234 => (x"ca",x"1e",x"49",x"69"),
  1235 => (x"c0",x"49",x"12",x"82"),
  1236 => (x"c0",x"87",x"e0",x"e6"),
  1237 => (x"87",x"c9",x"d4",x"49"),
  1238 => (x"f8",x"c0",x"49",x"74"),
  1239 => (x"8e",x"f8",x"87",x"e7"),
  1240 => (x"1e",x"87",x"f8",x"f4"),
  1241 => (x"4b",x"71",x"1e",x"73"),
  1242 => (x"87",x"c3",x"ff",x"49"),
  1243 => (x"fe",x"fe",x"49",x"73"),
  1244 => (x"87",x"e9",x"f4",x"87"),
  1245 => (x"71",x"1e",x"73",x"1e"),
  1246 => (x"4a",x"a3",x"c6",x"4b"),
  1247 => (x"c1",x"87",x"db",x"02"),
  1248 => (x"87",x"d6",x"02",x"8a"),
  1249 => (x"da",x"c1",x"02",x"8a"),
  1250 => (x"c0",x"02",x"8a",x"87"),
  1251 => (x"02",x"8a",x"87",x"fc"),
  1252 => (x"8a",x"87",x"e1",x"c0"),
  1253 => (x"c1",x"87",x"cb",x"02"),
  1254 => (x"49",x"c7",x"87",x"db"),
  1255 => (x"c1",x"87",x"c0",x"fd"),
  1256 => (x"c5",x"c3",x"87",x"de"),
  1257 => (x"c1",x"02",x"bf",x"d0"),
  1258 => (x"c1",x"48",x"87",x"cb"),
  1259 => (x"d4",x"c5",x"c3",x"88"),
  1260 => (x"87",x"c1",x"c1",x"58"),
  1261 => (x"bf",x"d4",x"c5",x"c3"),
  1262 => (x"87",x"f9",x"c0",x"02"),
  1263 => (x"bf",x"d0",x"c5",x"c3"),
  1264 => (x"c3",x"80",x"c1",x"48"),
  1265 => (x"c0",x"58",x"d4",x"c5"),
  1266 => (x"c5",x"c3",x"87",x"eb"),
  1267 => (x"c6",x"49",x"bf",x"d0"),
  1268 => (x"d4",x"c5",x"c3",x"89"),
  1269 => (x"a9",x"b7",x"c0",x"59"),
  1270 => (x"c3",x"87",x"da",x"03"),
  1271 => (x"c0",x"48",x"d0",x"c5"),
  1272 => (x"c3",x"87",x"d2",x"78"),
  1273 => (x"02",x"bf",x"d4",x"c5"),
  1274 => (x"c5",x"c3",x"87",x"cb"),
  1275 => (x"c6",x"48",x"bf",x"d0"),
  1276 => (x"d4",x"c5",x"c3",x"80"),
  1277 => (x"d1",x"49",x"c0",x"58"),
  1278 => (x"49",x"73",x"87",x"e7"),
  1279 => (x"87",x"c5",x"f6",x"c0"),
  1280 => (x"0e",x"87",x"da",x"f2"),
  1281 => (x"0e",x"5c",x"5b",x"5e"),
  1282 => (x"66",x"cc",x"4c",x"71"),
  1283 => (x"cb",x"4b",x"74",x"1e"),
  1284 => (x"f7",x"e4",x"c1",x"93"),
  1285 => (x"4a",x"a3",x"c4",x"83"),
  1286 => (x"f2",x"fe",x"49",x"6a"),
  1287 => (x"ca",x"c1",x"87",x"da"),
  1288 => (x"a3",x"c8",x"7b",x"dd"),
  1289 => (x"51",x"66",x"d4",x"49"),
  1290 => (x"d8",x"49",x"a3",x"c9"),
  1291 => (x"a3",x"ca",x"51",x"66"),
  1292 => (x"51",x"66",x"dc",x"49"),
  1293 => (x"87",x"e3",x"f1",x"26"),
  1294 => (x"5c",x"5b",x"5e",x"0e"),
  1295 => (x"d0",x"ff",x"0e",x"5d"),
  1296 => (x"59",x"a6",x"d8",x"86"),
  1297 => (x"c0",x"48",x"a6",x"c4"),
  1298 => (x"c1",x"80",x"c4",x"78"),
  1299 => (x"c4",x"78",x"66",x"c4"),
  1300 => (x"c4",x"78",x"c1",x"80"),
  1301 => (x"c3",x"78",x"c1",x"80"),
  1302 => (x"c1",x"48",x"d4",x"c5"),
  1303 => (x"cc",x"c5",x"c3",x"78"),
  1304 => (x"a8",x"de",x"48",x"bf"),
  1305 => (x"f3",x"87",x"cb",x"05"),
  1306 => (x"49",x"70",x"87",x"e5"),
  1307 => (x"ce",x"59",x"a6",x"c8"),
  1308 => (x"ed",x"e8",x"87",x"f8"),
  1309 => (x"87",x"cf",x"e9",x"87"),
  1310 => (x"70",x"87",x"dc",x"e8"),
  1311 => (x"ac",x"fb",x"c0",x"4c"),
  1312 => (x"87",x"d0",x"c1",x"02"),
  1313 => (x"c1",x"05",x"66",x"d4"),
  1314 => (x"1e",x"c0",x"87",x"c2"),
  1315 => (x"c1",x"1e",x"c1",x"1e"),
  1316 => (x"c0",x"1e",x"da",x"e6"),
  1317 => (x"87",x"eb",x"fd",x"49"),
  1318 => (x"4a",x"66",x"d0",x"c1"),
  1319 => (x"49",x"6a",x"82",x"c4"),
  1320 => (x"51",x"74",x"81",x"c7"),
  1321 => (x"1e",x"d8",x"1e",x"c1"),
  1322 => (x"81",x"c8",x"49",x"6a"),
  1323 => (x"d8",x"87",x"ec",x"e8"),
  1324 => (x"66",x"c4",x"c1",x"86"),
  1325 => (x"01",x"a8",x"c0",x"48"),
  1326 => (x"a6",x"c4",x"87",x"c7"),
  1327 => (x"ce",x"78",x"c1",x"48"),
  1328 => (x"66",x"c4",x"c1",x"87"),
  1329 => (x"cc",x"88",x"c1",x"48"),
  1330 => (x"87",x"c3",x"58",x"a6"),
  1331 => (x"cc",x"87",x"f8",x"e7"),
  1332 => (x"78",x"c2",x"48",x"a6"),
  1333 => (x"cd",x"02",x"9c",x"74"),
  1334 => (x"66",x"c4",x"87",x"cc"),
  1335 => (x"66",x"c8",x"c1",x"48"),
  1336 => (x"c1",x"cd",x"03",x"a8"),
  1337 => (x"48",x"a6",x"d8",x"87"),
  1338 => (x"ea",x"e6",x"78",x"c0"),
  1339 => (x"c1",x"4c",x"70",x"87"),
  1340 => (x"c2",x"05",x"ac",x"d0"),
  1341 => (x"66",x"d8",x"87",x"d6"),
  1342 => (x"87",x"ce",x"e9",x"7e"),
  1343 => (x"a6",x"dc",x"49",x"70"),
  1344 => (x"87",x"d3",x"e6",x"59"),
  1345 => (x"ec",x"c0",x"4c",x"70"),
  1346 => (x"ea",x"c1",x"05",x"ac"),
  1347 => (x"49",x"66",x"c4",x"87"),
  1348 => (x"c0",x"c1",x"91",x"cb"),
  1349 => (x"a1",x"c4",x"81",x"66"),
  1350 => (x"c8",x"4d",x"6a",x"4a"),
  1351 => (x"66",x"d8",x"4a",x"a1"),
  1352 => (x"df",x"cb",x"c1",x"52"),
  1353 => (x"87",x"ef",x"e5",x"79"),
  1354 => (x"02",x"9c",x"4c",x"70"),
  1355 => (x"fb",x"c0",x"87",x"d8"),
  1356 => (x"87",x"d2",x"02",x"ac"),
  1357 => (x"de",x"e5",x"55",x"74"),
  1358 => (x"9c",x"4c",x"70",x"87"),
  1359 => (x"c0",x"87",x"c7",x"02"),
  1360 => (x"ff",x"05",x"ac",x"fb"),
  1361 => (x"e0",x"c0",x"87",x"ee"),
  1362 => (x"55",x"c1",x"c2",x"55"),
  1363 => (x"d4",x"7d",x"97",x"c0"),
  1364 => (x"a9",x"6e",x"49",x"66"),
  1365 => (x"c4",x"87",x"db",x"05"),
  1366 => (x"66",x"c8",x"48",x"66"),
  1367 => (x"87",x"ca",x"04",x"a8"),
  1368 => (x"c1",x"48",x"66",x"c4"),
  1369 => (x"58",x"a6",x"c8",x"80"),
  1370 => (x"66",x"c8",x"87",x"c8"),
  1371 => (x"cc",x"88",x"c1",x"48"),
  1372 => (x"e2",x"e4",x"58",x"a6"),
  1373 => (x"c1",x"4c",x"70",x"87"),
  1374 => (x"c8",x"05",x"ac",x"d0"),
  1375 => (x"48",x"66",x"d0",x"87"),
  1376 => (x"a6",x"d4",x"80",x"c1"),
  1377 => (x"ac",x"d0",x"c1",x"58"),
  1378 => (x"87",x"ea",x"fd",x"02"),
  1379 => (x"d4",x"48",x"a6",x"dc"),
  1380 => (x"66",x"d8",x"78",x"66"),
  1381 => (x"a8",x"66",x"dc",x"48"),
  1382 => (x"87",x"dc",x"c9",x"05"),
  1383 => (x"48",x"a6",x"e0",x"c0"),
  1384 => (x"c4",x"78",x"f0",x"c0"),
  1385 => (x"78",x"66",x"cc",x"80"),
  1386 => (x"78",x"c0",x"80",x"c4"),
  1387 => (x"c0",x"48",x"74",x"7e"),
  1388 => (x"f0",x"c0",x"88",x"fb"),
  1389 => (x"98",x"70",x"58",x"a6"),
  1390 => (x"87",x"d7",x"c8",x"02"),
  1391 => (x"c0",x"88",x"cb",x"48"),
  1392 => (x"70",x"58",x"a6",x"f0"),
  1393 => (x"e9",x"c0",x"02",x"98"),
  1394 => (x"88",x"c9",x"48",x"87"),
  1395 => (x"58",x"a6",x"f0",x"c0"),
  1396 => (x"c3",x"02",x"98",x"70"),
  1397 => (x"c4",x"48",x"87",x"e1"),
  1398 => (x"a6",x"f0",x"c0",x"88"),
  1399 => (x"02",x"98",x"70",x"58"),
  1400 => (x"c1",x"48",x"87",x"d6"),
  1401 => (x"a6",x"f0",x"c0",x"88"),
  1402 => (x"02",x"98",x"70",x"58"),
  1403 => (x"c7",x"87",x"c8",x"c3"),
  1404 => (x"e0",x"c0",x"87",x"db"),
  1405 => (x"78",x"c0",x"48",x"a6"),
  1406 => (x"c1",x"48",x"66",x"cc"),
  1407 => (x"58",x"a6",x"d0",x"80"),
  1408 => (x"70",x"87",x"d4",x"e2"),
  1409 => (x"ac",x"ec",x"c0",x"4c"),
  1410 => (x"c0",x"87",x"d5",x"02"),
  1411 => (x"c6",x"02",x"66",x"e0"),
  1412 => (x"a6",x"e4",x"c0",x"87"),
  1413 => (x"74",x"87",x"c9",x"5c"),
  1414 => (x"88",x"f0",x"c0",x"48"),
  1415 => (x"58",x"a6",x"e8",x"c0"),
  1416 => (x"02",x"ac",x"ec",x"c0"),
  1417 => (x"ee",x"e1",x"87",x"cc"),
  1418 => (x"c0",x"4c",x"70",x"87"),
  1419 => (x"ff",x"05",x"ac",x"ec"),
  1420 => (x"e0",x"c0",x"87",x"f4"),
  1421 => (x"66",x"d4",x"1e",x"66"),
  1422 => (x"ec",x"c0",x"1e",x"49"),
  1423 => (x"e6",x"c1",x"1e",x"66"),
  1424 => (x"66",x"d4",x"1e",x"da"),
  1425 => (x"87",x"fb",x"f6",x"49"),
  1426 => (x"1e",x"ca",x"1e",x"c0"),
  1427 => (x"cb",x"49",x"66",x"dc"),
  1428 => (x"66",x"d8",x"c1",x"91"),
  1429 => (x"48",x"a6",x"d8",x"81"),
  1430 => (x"d8",x"78",x"a1",x"c4"),
  1431 => (x"e1",x"49",x"bf",x"66"),
  1432 => (x"86",x"d8",x"87",x"f9"),
  1433 => (x"06",x"a8",x"b7",x"c0"),
  1434 => (x"c1",x"87",x"c7",x"c1"),
  1435 => (x"c8",x"1e",x"de",x"1e"),
  1436 => (x"e1",x"49",x"bf",x"66"),
  1437 => (x"86",x"c8",x"87",x"e5"),
  1438 => (x"c0",x"48",x"49",x"70"),
  1439 => (x"e4",x"c0",x"88",x"08"),
  1440 => (x"b7",x"c0",x"58",x"a6"),
  1441 => (x"e9",x"c0",x"06",x"a8"),
  1442 => (x"66",x"e0",x"c0",x"87"),
  1443 => (x"a8",x"b7",x"dd",x"48"),
  1444 => (x"6e",x"87",x"df",x"03"),
  1445 => (x"e0",x"c0",x"49",x"bf"),
  1446 => (x"e0",x"c0",x"81",x"66"),
  1447 => (x"c1",x"49",x"66",x"51"),
  1448 => (x"81",x"bf",x"6e",x"81"),
  1449 => (x"c0",x"51",x"c1",x"c2"),
  1450 => (x"c2",x"49",x"66",x"e0"),
  1451 => (x"81",x"bf",x"6e",x"81"),
  1452 => (x"7e",x"c1",x"51",x"c0"),
  1453 => (x"e2",x"87",x"dc",x"c4"),
  1454 => (x"e4",x"c0",x"87",x"d0"),
  1455 => (x"c9",x"e2",x"58",x"a6"),
  1456 => (x"a6",x"e8",x"c0",x"87"),
  1457 => (x"a8",x"ec",x"c0",x"58"),
  1458 => (x"87",x"cb",x"c0",x"05"),
  1459 => (x"48",x"a6",x"e4",x"c0"),
  1460 => (x"78",x"66",x"e0",x"c0"),
  1461 => (x"ff",x"87",x"c4",x"c0"),
  1462 => (x"c4",x"87",x"fc",x"de"),
  1463 => (x"91",x"cb",x"49",x"66"),
  1464 => (x"48",x"66",x"c0",x"c1"),
  1465 => (x"7e",x"70",x"80",x"71"),
  1466 => (x"82",x"c8",x"4a",x"6e"),
  1467 => (x"81",x"ca",x"49",x"6e"),
  1468 => (x"51",x"66",x"e0",x"c0"),
  1469 => (x"49",x"66",x"e4",x"c0"),
  1470 => (x"e0",x"c0",x"81",x"c1"),
  1471 => (x"48",x"c1",x"89",x"66"),
  1472 => (x"49",x"70",x"30",x"71"),
  1473 => (x"97",x"71",x"89",x"c1"),
  1474 => (x"c1",x"c9",x"c3",x"7a"),
  1475 => (x"e0",x"c0",x"49",x"bf"),
  1476 => (x"6a",x"97",x"29",x"66"),
  1477 => (x"98",x"71",x"48",x"4a"),
  1478 => (x"58",x"a6",x"f0",x"c0"),
  1479 => (x"81",x"c4",x"49",x"6e"),
  1480 => (x"66",x"dc",x"4d",x"69"),
  1481 => (x"a8",x"66",x"d8",x"48"),
  1482 => (x"87",x"c8",x"c0",x"02"),
  1483 => (x"c0",x"48",x"a6",x"d8"),
  1484 => (x"87",x"c5",x"c0",x"78"),
  1485 => (x"c1",x"48",x"a6",x"d8"),
  1486 => (x"1e",x"66",x"d8",x"78"),
  1487 => (x"75",x"1e",x"e0",x"c0"),
  1488 => (x"d6",x"de",x"ff",x"49"),
  1489 => (x"70",x"86",x"c8",x"87"),
  1490 => (x"ac",x"b7",x"c0",x"4c"),
  1491 => (x"87",x"d4",x"c1",x"06"),
  1492 => (x"e0",x"c0",x"85",x"74"),
  1493 => (x"75",x"89",x"74",x"49"),
  1494 => (x"de",x"e1",x"c1",x"4b"),
  1495 => (x"e5",x"fe",x"71",x"4a"),
  1496 => (x"85",x"c2",x"87",x"c6"),
  1497 => (x"48",x"66",x"e8",x"c0"),
  1498 => (x"ec",x"c0",x"80",x"c1"),
  1499 => (x"ec",x"c0",x"58",x"a6"),
  1500 => (x"81",x"c1",x"49",x"66"),
  1501 => (x"c0",x"02",x"a9",x"70"),
  1502 => (x"a6",x"d8",x"87",x"c8"),
  1503 => (x"c0",x"78",x"c0",x"48"),
  1504 => (x"a6",x"d8",x"87",x"c5"),
  1505 => (x"d8",x"78",x"c1",x"48"),
  1506 => (x"a4",x"c2",x"1e",x"66"),
  1507 => (x"48",x"e0",x"c0",x"49"),
  1508 => (x"49",x"70",x"88",x"71"),
  1509 => (x"ff",x"49",x"75",x"1e"),
  1510 => (x"c8",x"87",x"c0",x"dd"),
  1511 => (x"a8",x"b7",x"c0",x"86"),
  1512 => (x"87",x"c0",x"ff",x"01"),
  1513 => (x"02",x"66",x"e8",x"c0"),
  1514 => (x"6e",x"87",x"d1",x"c0"),
  1515 => (x"c0",x"81",x"c9",x"49"),
  1516 => (x"6e",x"51",x"66",x"e8"),
  1517 => (x"ef",x"cc",x"c1",x"48"),
  1518 => (x"87",x"cc",x"c0",x"78"),
  1519 => (x"81",x"c9",x"49",x"6e"),
  1520 => (x"48",x"6e",x"51",x"c2"),
  1521 => (x"78",x"e3",x"cd",x"c1"),
  1522 => (x"c6",x"c0",x"7e",x"c1"),
  1523 => (x"f6",x"db",x"ff",x"87"),
  1524 => (x"6e",x"4c",x"70",x"87"),
  1525 => (x"87",x"f5",x"c0",x"02"),
  1526 => (x"c8",x"48",x"66",x"c4"),
  1527 => (x"c0",x"04",x"a8",x"66"),
  1528 => (x"66",x"c4",x"87",x"cb"),
  1529 => (x"c8",x"80",x"c1",x"48"),
  1530 => (x"e0",x"c0",x"58",x"a6"),
  1531 => (x"48",x"66",x"c8",x"87"),
  1532 => (x"a6",x"cc",x"88",x"c1"),
  1533 => (x"87",x"d5",x"c0",x"58"),
  1534 => (x"05",x"ac",x"c6",x"c1"),
  1535 => (x"cc",x"87",x"c8",x"c0"),
  1536 => (x"80",x"c1",x"48",x"66"),
  1537 => (x"ff",x"58",x"a6",x"d0"),
  1538 => (x"70",x"87",x"fc",x"da"),
  1539 => (x"48",x"66",x"d0",x"4c"),
  1540 => (x"a6",x"d4",x"80",x"c1"),
  1541 => (x"02",x"9c",x"74",x"58"),
  1542 => (x"c4",x"87",x"cb",x"c0"),
  1543 => (x"c8",x"c1",x"48",x"66"),
  1544 => (x"f2",x"04",x"a8",x"66"),
  1545 => (x"da",x"ff",x"87",x"ff"),
  1546 => (x"66",x"c4",x"87",x"d4"),
  1547 => (x"03",x"a8",x"c7",x"48"),
  1548 => (x"c3",x"87",x"e5",x"c0"),
  1549 => (x"c0",x"48",x"d4",x"c5"),
  1550 => (x"49",x"66",x"c4",x"78"),
  1551 => (x"c0",x"c1",x"91",x"cb"),
  1552 => (x"a1",x"c4",x"81",x"66"),
  1553 => (x"c0",x"4a",x"6a",x"4a"),
  1554 => (x"66",x"c4",x"79",x"52"),
  1555 => (x"c8",x"80",x"c1",x"48"),
  1556 => (x"a8",x"c7",x"58",x"a6"),
  1557 => (x"87",x"db",x"ff",x"04"),
  1558 => (x"e0",x"8e",x"d0",x"ff"),
  1559 => (x"20",x"3a",x"87",x"fb"),
  1560 => (x"1e",x"73",x"1e",x"00"),
  1561 => (x"02",x"9b",x"4b",x"71"),
  1562 => (x"c5",x"c3",x"87",x"c6"),
  1563 => (x"78",x"c0",x"48",x"d0"),
  1564 => (x"c5",x"c3",x"1e",x"c7"),
  1565 => (x"1e",x"49",x"bf",x"d0"),
  1566 => (x"1e",x"f7",x"e4",x"c1"),
  1567 => (x"bf",x"cc",x"c5",x"c3"),
  1568 => (x"87",x"f4",x"ee",x"49"),
  1569 => (x"c5",x"c3",x"86",x"cc"),
  1570 => (x"e9",x"49",x"bf",x"cc"),
  1571 => (x"9b",x"73",x"87",x"f9"),
  1572 => (x"c1",x"87",x"c8",x"02"),
  1573 => (x"c0",x"49",x"f7",x"e4"),
  1574 => (x"ff",x"87",x"fc",x"e4"),
  1575 => (x"1e",x"87",x"fe",x"df"),
  1576 => (x"c1",x"87",x"d6",x"c7"),
  1577 => (x"87",x"f9",x"fe",x"49"),
  1578 => (x"87",x"f4",x"e9",x"fe"),
  1579 => (x"cd",x"02",x"98",x"70"),
  1580 => (x"f1",x"f2",x"fe",x"87"),
  1581 => (x"02",x"98",x"70",x"87"),
  1582 => (x"4a",x"c1",x"87",x"c4"),
  1583 => (x"4a",x"c0",x"87",x"c2"),
  1584 => (x"ce",x"05",x"9a",x"72"),
  1585 => (x"c1",x"1e",x"c0",x"87"),
  1586 => (x"c0",x"49",x"f0",x"e3"),
  1587 => (x"c4",x"87",x"ff",x"f2"),
  1588 => (x"c0",x"87",x"fe",x"86"),
  1589 => (x"fb",x"e3",x"c1",x"1e"),
  1590 => (x"f1",x"f2",x"c0",x"49"),
  1591 => (x"c1",x"1e",x"c0",x"87"),
  1592 => (x"70",x"87",x"c8",x"cf"),
  1593 => (x"e5",x"f2",x"c0",x"49"),
  1594 => (x"87",x"cc",x"c3",x"87"),
  1595 => (x"4f",x"26",x"8e",x"f8"),
  1596 => (x"66",x"20",x"44",x"53"),
  1597 => (x"65",x"6c",x"69",x"61"),
  1598 => (x"42",x"00",x"2e",x"64"),
  1599 => (x"69",x"74",x"6f",x"6f"),
  1600 => (x"2e",x"2e",x"67",x"6e"),
  1601 => (x"c0",x"1e",x"00",x"2e"),
  1602 => (x"c0",x"87",x"f0",x"e7"),
  1603 => (x"f6",x"87",x"ca",x"f6"),
  1604 => (x"1e",x"4f",x"26",x"87"),
  1605 => (x"48",x"d0",x"c5",x"c3"),
  1606 => (x"c5",x"c3",x"78",x"c0"),
  1607 => (x"78",x"c0",x"48",x"cc"),
  1608 => (x"e1",x"87",x"fc",x"fd"),
  1609 => (x"26",x"48",x"c0",x"87"),
  1610 => (x"45",x"20",x"80",x"4f"),
  1611 => (x"00",x"74",x"69",x"78"),
  1612 => (x"61",x"42",x"20",x"80"),
  1613 => (x"df",x"00",x"6b",x"63"),
  1614 => (x"65",x"00",x"00",x"12"),
  1615 => (x"00",x"00",x"00",x"31"),
  1616 => (x"12",x"df",x"00",x"00"),
  1617 => (x"31",x"83",x"00",x"00"),
  1618 => (x"00",x"00",x"00",x"00"),
  1619 => (x"00",x"12",x"df",x"00"),
  1620 => (x"00",x"31",x"a1",x"00"),
  1621 => (x"00",x"00",x"00",x"00"),
  1622 => (x"00",x"00",x"12",x"df"),
  1623 => (x"00",x"00",x"31",x"bf"),
  1624 => (x"df",x"00",x"00",x"00"),
  1625 => (x"dd",x"00",x"00",x"12"),
  1626 => (x"00",x"00",x"00",x"31"),
  1627 => (x"12",x"df",x"00",x"00"),
  1628 => (x"31",x"fb",x"00",x"00"),
  1629 => (x"00",x"00",x"00",x"00"),
  1630 => (x"00",x"12",x"df",x"00"),
  1631 => (x"00",x"32",x"19",x"00"),
  1632 => (x"00",x"00",x"00",x"00"),
  1633 => (x"00",x"00",x"12",x"df"),
  1634 => (x"00",x"00",x"00",x"00"),
  1635 => (x"74",x"00",x"00",x"00"),
  1636 => (x"00",x"00",x"00",x"13"),
  1637 => (x"00",x"00",x"00",x"00"),
  1638 => (x"6f",x"4c",x"00",x"00"),
  1639 => (x"2a",x"20",x"64",x"61"),
  1640 => (x"fe",x"1e",x"00",x"2e"),
  1641 => (x"78",x"c0",x"48",x"f0"),
  1642 => (x"09",x"79",x"09",x"cd"),
  1643 => (x"1e",x"1e",x"4f",x"26"),
  1644 => (x"7e",x"bf",x"f0",x"fe"),
  1645 => (x"4f",x"26",x"26",x"48"),
  1646 => (x"48",x"f0",x"fe",x"1e"),
  1647 => (x"4f",x"26",x"78",x"c1"),
  1648 => (x"48",x"f0",x"fe",x"1e"),
  1649 => (x"4f",x"26",x"78",x"c0"),
  1650 => (x"c0",x"4a",x"71",x"1e"),
  1651 => (x"4f",x"26",x"52",x"52"),
  1652 => (x"5c",x"5b",x"5e",x"0e"),
  1653 => (x"86",x"f4",x"0e",x"5d"),
  1654 => (x"6d",x"97",x"4d",x"71"),
  1655 => (x"4c",x"a5",x"c1",x"7e"),
  1656 => (x"c8",x"48",x"6c",x"97"),
  1657 => (x"48",x"6e",x"58",x"a6"),
  1658 => (x"05",x"a8",x"66",x"c4"),
  1659 => (x"48",x"ff",x"87",x"c5"),
  1660 => (x"ff",x"87",x"e6",x"c0"),
  1661 => (x"a5",x"c2",x"87",x"ca"),
  1662 => (x"4b",x"6c",x"97",x"49"),
  1663 => (x"97",x"4b",x"a3",x"71"),
  1664 => (x"6c",x"97",x"4b",x"6b"),
  1665 => (x"c1",x"48",x"6e",x"7e"),
  1666 => (x"58",x"a6",x"c8",x"80"),
  1667 => (x"a6",x"cc",x"98",x"c7"),
  1668 => (x"7c",x"97",x"70",x"58"),
  1669 => (x"73",x"87",x"e1",x"fe"),
  1670 => (x"26",x"8e",x"f4",x"48"),
  1671 => (x"26",x"4c",x"26",x"4d"),
  1672 => (x"0e",x"4f",x"26",x"4b"),
  1673 => (x"0e",x"5c",x"5b",x"5e"),
  1674 => (x"4c",x"71",x"86",x"f4"),
  1675 => (x"c3",x"4a",x"66",x"d8"),
  1676 => (x"a4",x"c2",x"9a",x"ff"),
  1677 => (x"49",x"6c",x"97",x"4b"),
  1678 => (x"72",x"49",x"a1",x"73"),
  1679 => (x"7e",x"6c",x"97",x"51"),
  1680 => (x"80",x"c1",x"48",x"6e"),
  1681 => (x"c7",x"58",x"a6",x"c8"),
  1682 => (x"58",x"a6",x"cc",x"98"),
  1683 => (x"8e",x"f4",x"54",x"70"),
  1684 => (x"1e",x"87",x"ca",x"ff"),
  1685 => (x"87",x"e8",x"fd",x"1e"),
  1686 => (x"49",x"4a",x"bf",x"e0"),
  1687 => (x"99",x"c0",x"e0",x"c0"),
  1688 => (x"72",x"87",x"cb",x"02"),
  1689 => (x"f7",x"c8",x"c3",x"1e"),
  1690 => (x"87",x"f7",x"fe",x"49"),
  1691 => (x"fd",x"fc",x"86",x"c4"),
  1692 => (x"fd",x"7e",x"70",x"87"),
  1693 => (x"26",x"26",x"87",x"c2"),
  1694 => (x"c8",x"c3",x"1e",x"4f"),
  1695 => (x"c7",x"fd",x"49",x"f7"),
  1696 => (x"d3",x"e9",x"c1",x"87"),
  1697 => (x"87",x"da",x"fc",x"49"),
  1698 => (x"26",x"87",x"d0",x"c5"),
  1699 => (x"5b",x"5e",x"0e",x"4f"),
  1700 => (x"c3",x"0e",x"5d",x"5c"),
  1701 => (x"4a",x"bf",x"d6",x"c9"),
  1702 => (x"bf",x"e1",x"eb",x"c1"),
  1703 => (x"bc",x"72",x"4c",x"49"),
  1704 => (x"db",x"fc",x"4d",x"71"),
  1705 => (x"74",x"4b",x"c0",x"87"),
  1706 => (x"02",x"99",x"d0",x"49"),
  1707 => (x"49",x"75",x"87",x"d5"),
  1708 => (x"1e",x"71",x"99",x"d0"),
  1709 => (x"f1",x"c1",x"1e",x"c0"),
  1710 => (x"82",x"73",x"4a",x"ea"),
  1711 => (x"e4",x"c0",x"49",x"12"),
  1712 => (x"c1",x"86",x"c8",x"87"),
  1713 => (x"c8",x"83",x"2d",x"2c"),
  1714 => (x"da",x"ff",x"04",x"ab"),
  1715 => (x"87",x"e8",x"fb",x"87"),
  1716 => (x"48",x"e1",x"eb",x"c1"),
  1717 => (x"bf",x"d6",x"c9",x"c3"),
  1718 => (x"26",x"4d",x"26",x"78"),
  1719 => (x"26",x"4b",x"26",x"4c"),
  1720 => (x"00",x"00",x"00",x"4f"),
  1721 => (x"d0",x"ff",x"1e",x"00"),
  1722 => (x"78",x"e1",x"c8",x"48"),
  1723 => (x"c5",x"48",x"d4",x"ff"),
  1724 => (x"02",x"66",x"c4",x"78"),
  1725 => (x"e0",x"c3",x"87",x"c3"),
  1726 => (x"02",x"66",x"c8",x"78"),
  1727 => (x"d4",x"ff",x"87",x"c6"),
  1728 => (x"78",x"f0",x"c3",x"48"),
  1729 => (x"71",x"48",x"d4",x"ff"),
  1730 => (x"48",x"d0",x"ff",x"78"),
  1731 => (x"c0",x"78",x"e1",x"c8"),
  1732 => (x"4f",x"26",x"78",x"e0"),
  1733 => (x"5c",x"5b",x"5e",x"0e"),
  1734 => (x"c3",x"4c",x"71",x"0e"),
  1735 => (x"fa",x"49",x"f7",x"c8"),
  1736 => (x"4a",x"70",x"87",x"ee"),
  1737 => (x"04",x"aa",x"b7",x"c0"),
  1738 => (x"c3",x"87",x"e3",x"c2"),
  1739 => (x"c9",x"05",x"aa",x"e0"),
  1740 => (x"d7",x"ef",x"c1",x"87"),
  1741 => (x"c2",x"78",x"c1",x"48"),
  1742 => (x"f0",x"c3",x"87",x"d4"),
  1743 => (x"87",x"c9",x"05",x"aa"),
  1744 => (x"48",x"d3",x"ef",x"c1"),
  1745 => (x"f5",x"c1",x"78",x"c1"),
  1746 => (x"d7",x"ef",x"c1",x"87"),
  1747 => (x"87",x"c7",x"02",x"bf"),
  1748 => (x"c0",x"c2",x"4b",x"72"),
  1749 => (x"72",x"87",x"c2",x"b3"),
  1750 => (x"05",x"9c",x"74",x"4b"),
  1751 => (x"ef",x"c1",x"87",x"d1"),
  1752 => (x"c1",x"1e",x"bf",x"d3"),
  1753 => (x"1e",x"bf",x"d7",x"ef"),
  1754 => (x"f8",x"fd",x"49",x"72"),
  1755 => (x"c1",x"86",x"c8",x"87"),
  1756 => (x"02",x"bf",x"d3",x"ef"),
  1757 => (x"73",x"87",x"e0",x"c0"),
  1758 => (x"29",x"b7",x"c4",x"49"),
  1759 => (x"ea",x"f0",x"c1",x"91"),
  1760 => (x"cf",x"4a",x"73",x"81"),
  1761 => (x"c1",x"92",x"c2",x"9a"),
  1762 => (x"70",x"30",x"72",x"48"),
  1763 => (x"72",x"ba",x"ff",x"4a"),
  1764 => (x"70",x"98",x"69",x"48"),
  1765 => (x"73",x"87",x"db",x"79"),
  1766 => (x"29",x"b7",x"c4",x"49"),
  1767 => (x"ea",x"f0",x"c1",x"91"),
  1768 => (x"cf",x"4a",x"73",x"81"),
  1769 => (x"c3",x"92",x"c2",x"9a"),
  1770 => (x"70",x"30",x"72",x"48"),
  1771 => (x"b0",x"69",x"48",x"4a"),
  1772 => (x"ef",x"c1",x"79",x"70"),
  1773 => (x"78",x"c0",x"48",x"d7"),
  1774 => (x"48",x"d3",x"ef",x"c1"),
  1775 => (x"c8",x"c3",x"78",x"c0"),
  1776 => (x"cb",x"f8",x"49",x"f7"),
  1777 => (x"c0",x"4a",x"70",x"87"),
  1778 => (x"fd",x"03",x"aa",x"b7"),
  1779 => (x"48",x"c0",x"87",x"dd"),
  1780 => (x"00",x"87",x"c8",x"fc"),
  1781 => (x"00",x"00",x"00",x"00"),
  1782 => (x"1e",x"00",x"00",x"00"),
  1783 => (x"49",x"72",x"4a",x"c0"),
  1784 => (x"f0",x"c1",x"91",x"c4"),
  1785 => (x"79",x"c0",x"81",x"ea"),
  1786 => (x"b7",x"d0",x"82",x"c1"),
  1787 => (x"87",x"ee",x"04",x"aa"),
  1788 => (x"5e",x"0e",x"4f",x"26"),
  1789 => (x"0e",x"5d",x"5c",x"5b"),
  1790 => (x"c3",x"f7",x"4d",x"71"),
  1791 => (x"c4",x"4a",x"75",x"87"),
  1792 => (x"c1",x"92",x"2a",x"b7"),
  1793 => (x"75",x"82",x"ea",x"f0"),
  1794 => (x"c2",x"9c",x"cf",x"4c"),
  1795 => (x"4b",x"49",x"6a",x"94"),
  1796 => (x"9b",x"c3",x"2b",x"74"),
  1797 => (x"30",x"74",x"48",x"c2"),
  1798 => (x"bc",x"ff",x"4c",x"70"),
  1799 => (x"98",x"71",x"48",x"74"),
  1800 => (x"d3",x"f6",x"7a",x"70"),
  1801 => (x"fa",x"48",x"73",x"87"),
  1802 => (x"00",x"00",x"87",x"ef"),
  1803 => (x"00",x"00",x"00",x"00"),
  1804 => (x"00",x"00",x"00",x"00"),
  1805 => (x"00",x"00",x"00",x"00"),
  1806 => (x"00",x"00",x"00",x"00"),
  1807 => (x"00",x"00",x"00",x"00"),
  1808 => (x"00",x"00",x"00",x"00"),
  1809 => (x"00",x"00",x"00",x"00"),
  1810 => (x"00",x"00",x"00",x"00"),
  1811 => (x"00",x"00",x"00",x"00"),
  1812 => (x"00",x"00",x"00",x"00"),
  1813 => (x"00",x"00",x"00",x"00"),
  1814 => (x"00",x"00",x"00",x"00"),
  1815 => (x"00",x"00",x"00",x"00"),
  1816 => (x"00",x"00",x"00",x"00"),
  1817 => (x"00",x"00",x"00",x"00"),
  1818 => (x"1e",x"16",x"00",x"00"),
  1819 => (x"36",x"2e",x"25",x"26"),
  1820 => (x"ff",x"1e",x"3e",x"3d"),
  1821 => (x"e1",x"c8",x"48",x"d0"),
  1822 => (x"ff",x"48",x"71",x"78"),
  1823 => (x"26",x"78",x"08",x"d4"),
  1824 => (x"d0",x"ff",x"1e",x"4f"),
  1825 => (x"78",x"e1",x"c8",x"48"),
  1826 => (x"d4",x"ff",x"48",x"71"),
  1827 => (x"66",x"c4",x"78",x"08"),
  1828 => (x"08",x"d4",x"ff",x"48"),
  1829 => (x"1e",x"4f",x"26",x"78"),
  1830 => (x"66",x"c4",x"4a",x"71"),
  1831 => (x"49",x"72",x"1e",x"49"),
  1832 => (x"ff",x"87",x"de",x"ff"),
  1833 => (x"e0",x"c0",x"48",x"d0"),
  1834 => (x"4f",x"26",x"26",x"78"),
  1835 => (x"c2",x"4a",x"71",x"1e"),
  1836 => (x"c3",x"03",x"aa",x"b7"),
  1837 => (x"87",x"c2",x"82",x"87"),
  1838 => (x"66",x"c4",x"82",x"ce"),
  1839 => (x"ff",x"49",x"72",x"1e"),
  1840 => (x"26",x"26",x"87",x"d5"),
  1841 => (x"d4",x"ff",x"1e",x"4f"),
  1842 => (x"7a",x"ff",x"c3",x"4a"),
  1843 => (x"c8",x"48",x"d0",x"ff"),
  1844 => (x"7a",x"de",x"78",x"e1"),
  1845 => (x"bf",x"c1",x"c9",x"c3"),
  1846 => (x"c8",x"48",x"49",x"7a"),
  1847 => (x"71",x"7a",x"70",x"28"),
  1848 => (x"70",x"28",x"d0",x"48"),
  1849 => (x"d8",x"48",x"71",x"7a"),
  1850 => (x"ff",x"7a",x"70",x"28"),
  1851 => (x"e0",x"c0",x"48",x"d0"),
  1852 => (x"0e",x"4f",x"26",x"78"),
  1853 => (x"5d",x"5c",x"5b",x"5e"),
  1854 => (x"c3",x"4c",x"71",x"0e"),
  1855 => (x"4d",x"bf",x"c1",x"c9"),
  1856 => (x"d0",x"2b",x"74",x"4b"),
  1857 => (x"83",x"c1",x"9b",x"66"),
  1858 => (x"04",x"ab",x"66",x"d4"),
  1859 => (x"4b",x"c0",x"87",x"c2"),
  1860 => (x"66",x"d0",x"4a",x"74"),
  1861 => (x"ff",x"31",x"72",x"49"),
  1862 => (x"73",x"99",x"75",x"b9"),
  1863 => (x"70",x"30",x"72",x"48"),
  1864 => (x"b0",x"71",x"48",x"4a"),
  1865 => (x"58",x"c5",x"c9",x"c3"),
  1866 => (x"26",x"87",x"da",x"fe"),
  1867 => (x"26",x"4c",x"26",x"4d"),
  1868 => (x"1e",x"4f",x"26",x"4b"),
  1869 => (x"c8",x"48",x"d0",x"ff"),
  1870 => (x"48",x"71",x"78",x"c9"),
  1871 => (x"78",x"08",x"d4",x"ff"),
  1872 => (x"71",x"1e",x"4f",x"26"),
  1873 => (x"87",x"eb",x"49",x"4a"),
  1874 => (x"c8",x"48",x"d0",x"ff"),
  1875 => (x"1e",x"4f",x"26",x"78"),
  1876 => (x"4b",x"71",x"1e",x"73"),
  1877 => (x"bf",x"d1",x"c9",x"c3"),
  1878 => (x"c2",x"87",x"c3",x"02"),
  1879 => (x"d0",x"ff",x"87",x"eb"),
  1880 => (x"78",x"c9",x"c8",x"48"),
  1881 => (x"e0",x"c0",x"49",x"73"),
  1882 => (x"48",x"d4",x"ff",x"b1"),
  1883 => (x"c9",x"c3",x"78",x"71"),
  1884 => (x"78",x"c0",x"48",x"c5"),
  1885 => (x"c5",x"02",x"66",x"c8"),
  1886 => (x"49",x"ff",x"c3",x"87"),
  1887 => (x"49",x"c0",x"87",x"c2"),
  1888 => (x"59",x"cd",x"c9",x"c3"),
  1889 => (x"c6",x"02",x"66",x"cc"),
  1890 => (x"d5",x"d5",x"c5",x"87"),
  1891 => (x"cf",x"87",x"c4",x"4a"),
  1892 => (x"c3",x"4a",x"ff",x"ff"),
  1893 => (x"c3",x"5a",x"d1",x"c9"),
  1894 => (x"c1",x"48",x"d1",x"c9"),
  1895 => (x"26",x"87",x"c4",x"78"),
  1896 => (x"26",x"4c",x"26",x"4d"),
  1897 => (x"0e",x"4f",x"26",x"4b"),
  1898 => (x"5d",x"5c",x"5b",x"5e"),
  1899 => (x"c3",x"4a",x"71",x"0e"),
  1900 => (x"4c",x"bf",x"cd",x"c9"),
  1901 => (x"cb",x"02",x"9a",x"72"),
  1902 => (x"91",x"c8",x"49",x"87"),
  1903 => (x"4b",x"c5",x"f5",x"c1"),
  1904 => (x"87",x"c4",x"83",x"71"),
  1905 => (x"4b",x"c5",x"f9",x"c1"),
  1906 => (x"49",x"13",x"4d",x"c0"),
  1907 => (x"c9",x"c3",x"99",x"74"),
  1908 => (x"ff",x"b9",x"bf",x"c9"),
  1909 => (x"78",x"71",x"48",x"d4"),
  1910 => (x"85",x"2c",x"b7",x"c1"),
  1911 => (x"04",x"ad",x"b7",x"c8"),
  1912 => (x"c9",x"c3",x"87",x"e8"),
  1913 => (x"c8",x"48",x"bf",x"c5"),
  1914 => (x"c9",x"c9",x"c3",x"80"),
  1915 => (x"87",x"ef",x"fe",x"58"),
  1916 => (x"71",x"1e",x"73",x"1e"),
  1917 => (x"9a",x"4a",x"13",x"4b"),
  1918 => (x"72",x"87",x"cb",x"02"),
  1919 => (x"87",x"e7",x"fe",x"49"),
  1920 => (x"05",x"9a",x"4a",x"13"),
  1921 => (x"da",x"fe",x"87",x"f5"),
  1922 => (x"c9",x"c3",x"1e",x"87"),
  1923 => (x"c3",x"49",x"bf",x"c5"),
  1924 => (x"c1",x"48",x"c5",x"c9"),
  1925 => (x"c0",x"c4",x"78",x"a1"),
  1926 => (x"db",x"03",x"a9",x"b7"),
  1927 => (x"48",x"d4",x"ff",x"87"),
  1928 => (x"bf",x"c9",x"c9",x"c3"),
  1929 => (x"c5",x"c9",x"c3",x"78"),
  1930 => (x"c9",x"c3",x"49",x"bf"),
  1931 => (x"a1",x"c1",x"48",x"c5"),
  1932 => (x"b7",x"c0",x"c4",x"78"),
  1933 => (x"87",x"e5",x"04",x"a9"),
  1934 => (x"c8",x"48",x"d0",x"ff"),
  1935 => (x"d1",x"c9",x"c3",x"78"),
  1936 => (x"26",x"78",x"c0",x"48"),
  1937 => (x"00",x"00",x"00",x"4f"),
  1938 => (x"00",x"00",x"00",x"00"),
  1939 => (x"00",x"00",x"00",x"00"),
  1940 => (x"00",x"00",x"5f",x"5f"),
  1941 => (x"03",x"03",x"00",x"00"),
  1942 => (x"00",x"03",x"03",x"00"),
  1943 => (x"7f",x"7f",x"14",x"00"),
  1944 => (x"14",x"7f",x"7f",x"14"),
  1945 => (x"2e",x"24",x"00",x"00"),
  1946 => (x"12",x"3a",x"6b",x"6b"),
  1947 => (x"36",x"6a",x"4c",x"00"),
  1948 => (x"32",x"56",x"6c",x"18"),
  1949 => (x"4f",x"7e",x"30",x"00"),
  1950 => (x"68",x"3a",x"77",x"59"),
  1951 => (x"04",x"00",x"00",x"40"),
  1952 => (x"00",x"00",x"03",x"07"),
  1953 => (x"1c",x"00",x"00",x"00"),
  1954 => (x"00",x"41",x"63",x"3e"),
  1955 => (x"41",x"00",x"00",x"00"),
  1956 => (x"00",x"1c",x"3e",x"63"),
  1957 => (x"3e",x"2a",x"08",x"00"),
  1958 => (x"2a",x"3e",x"1c",x"1c"),
  1959 => (x"08",x"08",x"00",x"08"),
  1960 => (x"08",x"08",x"3e",x"3e"),
  1961 => (x"80",x"00",x"00",x"00"),
  1962 => (x"00",x"00",x"60",x"e0"),
  1963 => (x"08",x"08",x"00",x"00"),
  1964 => (x"08",x"08",x"08",x"08"),
  1965 => (x"00",x"00",x"00",x"00"),
  1966 => (x"00",x"00",x"60",x"60"),
  1967 => (x"30",x"60",x"40",x"00"),
  1968 => (x"03",x"06",x"0c",x"18"),
  1969 => (x"7f",x"3e",x"00",x"01"),
  1970 => (x"3e",x"7f",x"4d",x"59"),
  1971 => (x"06",x"04",x"00",x"00"),
  1972 => (x"00",x"00",x"7f",x"7f"),
  1973 => (x"63",x"42",x"00",x"00"),
  1974 => (x"46",x"4f",x"59",x"71"),
  1975 => (x"63",x"22",x"00",x"00"),
  1976 => (x"36",x"7f",x"49",x"49"),
  1977 => (x"16",x"1c",x"18",x"00"),
  1978 => (x"10",x"7f",x"7f",x"13"),
  1979 => (x"67",x"27",x"00",x"00"),
  1980 => (x"39",x"7d",x"45",x"45"),
  1981 => (x"7e",x"3c",x"00",x"00"),
  1982 => (x"30",x"79",x"49",x"4b"),
  1983 => (x"01",x"01",x"00",x"00"),
  1984 => (x"07",x"0f",x"79",x"71"),
  1985 => (x"7f",x"36",x"00",x"00"),
  1986 => (x"36",x"7f",x"49",x"49"),
  1987 => (x"4f",x"06",x"00",x"00"),
  1988 => (x"1e",x"3f",x"69",x"49"),
  1989 => (x"00",x"00",x"00",x"00"),
  1990 => (x"00",x"00",x"66",x"66"),
  1991 => (x"80",x"00",x"00",x"00"),
  1992 => (x"00",x"00",x"66",x"e6"),
  1993 => (x"08",x"08",x"00",x"00"),
  1994 => (x"22",x"22",x"14",x"14"),
  1995 => (x"14",x"14",x"00",x"00"),
  1996 => (x"14",x"14",x"14",x"14"),
  1997 => (x"22",x"22",x"00",x"00"),
  1998 => (x"08",x"08",x"14",x"14"),
  1999 => (x"03",x"02",x"00",x"00"),
  2000 => (x"06",x"0f",x"59",x"51"),
  2001 => (x"41",x"7f",x"3e",x"00"),
  2002 => (x"1e",x"1f",x"55",x"5d"),
  2003 => (x"7f",x"7e",x"00",x"00"),
  2004 => (x"7e",x"7f",x"09",x"09"),
  2005 => (x"7f",x"7f",x"00",x"00"),
  2006 => (x"36",x"7f",x"49",x"49"),
  2007 => (x"3e",x"1c",x"00",x"00"),
  2008 => (x"41",x"41",x"41",x"63"),
  2009 => (x"7f",x"7f",x"00",x"00"),
  2010 => (x"1c",x"3e",x"63",x"41"),
  2011 => (x"7f",x"7f",x"00",x"00"),
  2012 => (x"41",x"41",x"49",x"49"),
  2013 => (x"7f",x"7f",x"00",x"00"),
  2014 => (x"01",x"01",x"09",x"09"),
  2015 => (x"7f",x"3e",x"00",x"00"),
  2016 => (x"7a",x"7b",x"49",x"41"),
  2017 => (x"7f",x"7f",x"00",x"00"),
  2018 => (x"7f",x"7f",x"08",x"08"),
  2019 => (x"41",x"00",x"00",x"00"),
  2020 => (x"00",x"41",x"7f",x"7f"),
  2021 => (x"60",x"20",x"00",x"00"),
  2022 => (x"3f",x"7f",x"40",x"40"),
  2023 => (x"08",x"7f",x"7f",x"00"),
  2024 => (x"41",x"63",x"36",x"1c"),
  2025 => (x"7f",x"7f",x"00",x"00"),
  2026 => (x"40",x"40",x"40",x"40"),
  2027 => (x"06",x"7f",x"7f",x"00"),
  2028 => (x"7f",x"7f",x"06",x"0c"),
  2029 => (x"06",x"7f",x"7f",x"00"),
  2030 => (x"7f",x"7f",x"18",x"0c"),
  2031 => (x"7f",x"3e",x"00",x"00"),
  2032 => (x"3e",x"7f",x"41",x"41"),
  2033 => (x"7f",x"7f",x"00",x"00"),
  2034 => (x"06",x"0f",x"09",x"09"),
  2035 => (x"41",x"7f",x"3e",x"00"),
  2036 => (x"40",x"7e",x"7f",x"61"),
  2037 => (x"7f",x"7f",x"00",x"00"),
  2038 => (x"66",x"7f",x"19",x"09"),
  2039 => (x"6f",x"26",x"00",x"00"),
  2040 => (x"32",x"7b",x"59",x"4d"),
  2041 => (x"01",x"01",x"00",x"00"),
  2042 => (x"01",x"01",x"7f",x"7f"),
  2043 => (x"7f",x"3f",x"00",x"00"),
  2044 => (x"3f",x"7f",x"40",x"40"),
  2045 => (x"3f",x"0f",x"00",x"00"),
  2046 => (x"0f",x"3f",x"70",x"70"),
  2047 => (x"30",x"7f",x"7f",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

